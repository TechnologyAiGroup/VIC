module s13207(CLK, SI, SE, g43, g49, g633, g634, g635, g645, g647, g648, g690, g694, g698, g702, g722, g723, g751, g752, g753, g754, g755, g756, g757, g781, g941, g962, g1000, g1008, g1016, g1080, g1234, g1553, g1554, SO, g206, g291, g372, g453, g534, g594, g785, g1006, g1015, g1017, g1246, g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829, g1870, g1871, g1894, g1911, g1944, g2662, g2844, g2888, g3077, g3096, g3130, g3159, g3191, g3829, g3859, g3860, g4267, g4316, g4370, g4371, g4372, g4373, g4655, g4657, g4660, g4661, g4663, g4664, g5143, g5164, g5571, g5669, g5678, g5682, g5684, g5687, g5729, g6207, g6212, g6223, g6236, g6269, g6425, g6648, g6653, g6675, g6849, g6850, g6895, g6909, g7048, g7063, g7103, g7283, g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291, g7292, g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504, g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732, g8216, g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958, g9128, g9132, g9204, g9280, g9297, g9299, g9305, g9308, g9310, g9312, g9314, g9378);
input CLK;
input SI;
input SE;
input g43;
input g49;
input g633;
input g634;
input g635;
input g645;
input g647;
input g648;
input g690;
input g694;
input g698;
input g702;
input g722;
input g723;
input g751;
input g752;
input g753;
input g754;
input g755;
input g756;
input g757;
input g781;
input g941;
input g962;
input g1000;
input g1008;
input g1016;
input g1080;
input g1234;
input g1553;
input g1554;
output SO;
output g206;
output g291;
output g372;
output g453;
output g534;
output g594;
output g785;
output g1006;
output g1015;
output g1017;
output g1246;
output g1724;
output g1783;
output g1798;
output g1804;
output g1810;
output g1817;
output g1824;
output g1829;
output g1870;
output g1871;
output g1894;
output g1911;
output g1944;
output g2662;
output g2844;
output g2888;
output g3077;
output g3096;
output g3130;
output g3159;
output g3191;
output g3829;
output g3859;
output g3860;
output g4267;
output g4316;
output g4370;
output g4371;
output g4372;
output g4373;
output g4655;
output g4657;
output g4660;
output g4661;
output g4663;
output g4664;
output g5143;
output g5164;
output g5571;
output g5669;
output g5678;
output g5682;
output g5684;
output g5687;
output g5729;
output g6207;
output g6212;
output g6223;
output g6236;
output g6269;
output g6425;
output g6648;
output g6653;
output g6675;
output g6849;
output g6850;
output g6895;
output g6909;
output g7048;
output g7063;
output g7103;
output g7283;
output g7284;
output g7285;
output g7286;
output g7287;
output g7288;
output g7289;
output g7290;
output g7291;
output g7292;
output g7293;
output g7294;
output g7295;
output g7298;
output g7423;
output g7424;
output g7425;
output g7474;
output g7504;
output g7505;
output g7506;
output g7507;
output g7508;
output g7514;
output g7729;
output g7730;
output g7731;
output g7732;
output g8216;
output g8217;
output g8218;
output g8219;
output g8234;
output g8661;
output g8663;
output g8872;
output g8958;
output g9128;
output g9132;
output g9204;
output g9280;
output g9297;
output g9299;
output g9305;
output g9308;
output g9310;
output g9312;
output g9314;
output g9378;
MUX2_X1 g_tmp_wire_0 (g6302, SI, SE, tmp_wire_0);
DFF_X1 g_g31 (tmp_wire_0, CLK, g31);
MUX2_X1 g_tmp_wire_1 (g6301, g31, SE, tmp_wire_1);
DFF_X1 g_g30 (tmp_wire_1, CLK, g30);
MUX2_X1 g_tmp_wire_2 (g6300, g30, SE, tmp_wire_2);
DFF_X1 g_g29 (tmp_wire_2, CLK, g29);
MUX2_X1 g_tmp_wire_3 (g6298, g29, SE, tmp_wire_3);
DFF_X1 g_g28 (tmp_wire_3, CLK, g28);
MUX2_X1 g_tmp_wire_4 (g6297, g28, SE, tmp_wire_4);
DFF_X1 g_g27 (tmp_wire_4, CLK, g27);
MUX2_X1 g_tmp_wire_5 (g6296, g27, SE, tmp_wire_5);
DFF_X1 g_g26 (tmp_wire_5, CLK, g26);
MUX2_X1 g_tmp_wire_6 (g6295, g26, SE, tmp_wire_6);
DFF_X1 g_g25 (tmp_wire_6, CLK, g25);
MUX2_X1 g_tmp_wire_7 (g6294, g25, SE, tmp_wire_7);
DFF_X1 g_g24 (tmp_wire_7, CLK, g24);
MUX2_X1 g_tmp_wire_8 (g6293, g24, SE, tmp_wire_8);
DFF_X1 g_g23 (tmp_wire_8, CLK, g23);
MUX2_X1 g_tmp_wire_9 (g6292, g23, SE, tmp_wire_9);
DFF_X1 g_g22 (tmp_wire_9, CLK, g22);
MUX2_X1 g_tmp_wire_10 (g8662, g22, SE, tmp_wire_10);
DFF_X1 g_g12 (tmp_wire_10, CLK, g12);
MUX2_X1 g_tmp_wire_11 (g6290, g12, SE, tmp_wire_11);
DFF_X1 g_g11 (tmp_wire_11, CLK, g11);
MUX2_X1 g_tmp_wire_12 (g6288, g11, SE, tmp_wire_12);
DFF_X1 g_g9 (tmp_wire_12, CLK, g9);
MUX2_X1 g_tmp_wire_13 (g9376, g9, SE, tmp_wire_13);
DFF_X1 g_g8 (tmp_wire_13, CLK, g8);
MUX2_X1 g_tmp_wire_14 (g9375, g8, SE, tmp_wire_14);
DFF_X1 g_g7 (tmp_wire_14, CLK, g7);
MUX2_X1 g_tmp_wire_15 (g9374, g7, SE, tmp_wire_15);
DFF_X1 g_g6 (tmp_wire_15, CLK, g6);
MUX2_X1 g_tmp_wire_16 (g9373, g6, SE, tmp_wire_16);
DFF_X1 g_g5 (tmp_wire_16, CLK, g5);
MUX2_X1 g_tmp_wire_17 (g9372, g5, SE, tmp_wire_17);
DFF_X1 g_g4 (tmp_wire_17, CLK, g4);
MUX2_X1 g_tmp_wire_18 (g9361, g4, SE, tmp_wire_18);
DFF_X1 g_g2 (tmp_wire_18, CLK, g2);
MUX2_X1 g_tmp_wire_19 (g9360, g2, SE, tmp_wire_19);
DFF_X1 g_g3 (tmp_wire_19, CLK, g3);
MUX2_X1 g_tmp_wire_20 (g9362, g3, SE, tmp_wire_20);
DFF_X1 g_g48 (tmp_wire_20, CLK, g48);
MUX2_X1 g_tmp_wire_21 (g6299, g48, SE, tmp_wire_21);
DFF_X1 g_g21 (tmp_wire_21, CLK, g21);
MUX2_X1 g_tmp_wire_22 (g6291, g21, SE, tmp_wire_22);
DFF_X1 g_g10 (tmp_wire_22, CLK, g10);
MUX2_X1 g_tmp_wire_23 (g6289, g10, SE, tmp_wire_23);
DFF_X1 g_g1 (tmp_wire_23, CLK, g1);
MUX2_X1 g_tmp_wire_24 (g9389, g1, SE, tmp_wire_24);
DFF_X1 g_g47 (tmp_wire_24, CLK, g47);
MUX2_X1 g_tmp_wire_25 (g8955, g47, SE, tmp_wire_25);
DFF_X1 g_g46 (tmp_wire_25, CLK, g46);
MUX2_X1 g_tmp_wire_26 (g6308, g46, SE, tmp_wire_26);
DFF_X1 g_g45 (tmp_wire_26, CLK, g45);
MUX2_X1 g_tmp_wire_27 (g6307, g45, SE, tmp_wire_27);
DFF_X1 g_g44 (tmp_wire_27, CLK, g44);
MUX2_X1 g_tmp_wire_28 (g6306, g44, SE, tmp_wire_28);
DFF_X1 g_g42 (tmp_wire_28, CLK, g42);
MUX2_X1 g_tmp_wire_29 (g6305, g42, SE, tmp_wire_29);
DFF_X1 g_g41 (tmp_wire_29, CLK, g41);
MUX2_X1 g_tmp_wire_30 (g6304, g41, SE, tmp_wire_30);
DFF_X1 g_g37 (tmp_wire_30, CLK, g37);
MUX2_X1 g_tmp_wire_31 (g6303, g37, SE, tmp_wire_31);
DFF_X1 g_g32 (tmp_wire_31, CLK, g32);
MUX2_X1 g_tmp_wire_32 (g5173, g32, SE, tmp_wire_32);
DFF_X1 g_g1207 (tmp_wire_32, CLK, g1207);
MUX2_X1 g_tmp_wire_33 (g5174, g1207, SE, tmp_wire_33);
DFF_X1 g_g1211 (tmp_wire_33, CLK, g1211);
MUX2_X1 g_tmp_wire_34 (g5736, g1211, SE, tmp_wire_34);
DFF_X1 g_g1214 (tmp_wire_34, CLK, g1214);
MUX2_X1 g_tmp_wire_35 (g6377, g1214, SE, tmp_wire_35);
DFF_X1 g_g1217 (tmp_wire_35, CLK, g1217);
MUX2_X1 g_tmp_wire_36 (g6378, g1217, SE, tmp_wire_36);
DFF_X1 g_g1220 (tmp_wire_36, CLK, g1220);
MUX2_X1 g_tmp_wire_37 (g6379, g1220, SE, tmp_wire_37);
DFF_X1 g_g1223 (tmp_wire_37, CLK, g1223);
MUX2_X1 g_tmp_wire_38 (g6857, g1223, SE, tmp_wire_38);
DFF_X1 g_g1224 (tmp_wire_38, CLK, g1224);
MUX2_X1 g_tmp_wire_39 (g6858, g1224, SE, tmp_wire_39);
DFF_X1 g_g1225 (tmp_wire_39, CLK, g1225);
MUX2_X1 g_tmp_wire_40 (g6859, g1225, SE, tmp_wire_40);
DFF_X1 g_g1226 (tmp_wire_40, CLK, g1226);
MUX2_X1 g_tmp_wire_41 (g7108, g1226, SE, tmp_wire_41);
DFF_X1 g_g1227 (tmp_wire_41, CLK, g1227);
MUX2_X1 g_tmp_wire_42 (g7109, g1227, SE, tmp_wire_42);
DFF_X1 g_g1228 (tmp_wire_42, CLK, g1228);
MUX2_X1 g_tmp_wire_43 (g7110, g1228, SE, tmp_wire_43);
DFF_X1 g_g1229 (tmp_wire_43, CLK, g1229);
MUX2_X1 g_tmp_wire_44 (g7300, g1229, SE, tmp_wire_44);
DFF_X1 g_g1230 (tmp_wire_44, CLK, g1230);
MUX2_X1 g_tmp_wire_45 (g1235, g1230, SE, tmp_wire_45);
DFF_X1 g_g1240 (tmp_wire_45, CLK, g1240);
MUX2_X1 g_tmp_wire_46 (g1240, g1240, SE, tmp_wire_46);
DFF_X1 g_g1236 (tmp_wire_46, CLK, g1236);
MUX2_X1 g_tmp_wire_47 (g1236, g1236, SE, tmp_wire_47);
DFF_X1 g_g1231 (tmp_wire_47, CLK, g1231);
MUX2_X1 g_tmp_wire_48 (g2659, g1231, SE, tmp_wire_48);
DFF_X1 g_g1244 (tmp_wire_48, CLK, g1244);
MUX2_X1 g_tmp_wire_49 (g1244, g1244, SE, tmp_wire_49);
DFF_X1 g_g1245 (tmp_wire_49, CLK, g1245);
MUX2_X1 g_tmp_wire_50 (g2660, g1245, SE, tmp_wire_50);
DFF_X1 g_g1243 (tmp_wire_50, CLK, g1243);
MUX2_X1 g_tmp_wire_51 (g6383, g1243, SE, tmp_wire_51);
DFF_X1 g_g1272 (tmp_wire_51, CLK, g1272);
MUX2_X1 g_tmp_wire_52 (g6384, g1272, SE, tmp_wire_52);
DFF_X1 g_g1276 (tmp_wire_52, CLK, g1276);
MUX2_X1 g_tmp_wire_53 (g7112, g1276, SE, tmp_wire_53);
DFF_X1 g_g1280 (tmp_wire_53, CLK, g1280);
MUX2_X1 g_tmp_wire_54 (g7301, g1280, SE, tmp_wire_54);
DFF_X1 g_g1284 (tmp_wire_54, CLK, g1284);
MUX2_X1 g_tmp_wire_55 (g7527, g1284, SE, tmp_wire_55);
DFF_X1 g_g1288 (tmp_wire_55, CLK, g1288);
MUX2_X1 g_tmp_wire_56 (g7302, g1288, SE, tmp_wire_56);
DFF_X1 g_g1292 (tmp_wire_56, CLK, g1292);
MUX2_X1 g_tmp_wire_57 (g7303, g1292, SE, tmp_wire_57);
DFF_X1 g_g1300 (tmp_wire_57, CLK, g1300);
MUX2_X1 g_tmp_wire_58 (g7304, g1300, SE, tmp_wire_58);
DFF_X1 g_g1296 (tmp_wire_58, CLK, g1296);
MUX2_X1 g_tmp_wire_59 (g5741, g1296, SE, tmp_wire_59);
DFF_X1 g_g1253 (tmp_wire_59, CLK, g1253);
MUX2_X1 g_tmp_wire_60 (g6385, g1253, SE, tmp_wire_60);
DFF_X1 g_g1308 (tmp_wire_60, CLK, g1308);
MUX2_X1 g_tmp_wire_61 (g1308, g1308, SE, tmp_wire_61);
DFF_X1 g_g1309 (tmp_wire_61, CLK, g1309);
MUX2_X1 g_tmp_wire_62 (g1309, g1309, SE, tmp_wire_62);
DFF_X1 g_g1310 (tmp_wire_62, CLK, g1310);
MUX2_X1 g_tmp_wire_63 (g1310, g1310, SE, tmp_wire_63);
DFF_X1 g_g1311 (tmp_wire_63, CLK, g1311);
MUX2_X1 g_tmp_wire_64 (g1311, g1311, SE, tmp_wire_64);
DFF_X1 g_g1312 (tmp_wire_64, CLK, g1312);
MUX2_X1 g_tmp_wire_65 (g1312, g1312, SE, tmp_wire_65);
DFF_X1 g_g1304 (tmp_wire_65, CLK, g1304);
MUX2_X1 g_tmp_wire_66 (g3858, g1304, SE, tmp_wire_66);
DFF_X1 g_g1307 (tmp_wire_66, CLK, g1307);
MUX2_X1 g_tmp_wire_67 (g6862, g1307, SE, tmp_wire_67);
DFF_X1 g_g1330 (tmp_wire_67, CLK, g1330);
MUX2_X1 g_tmp_wire_68 (g6863, g1330, SE, tmp_wire_68);
DFF_X1 g_g1333 (tmp_wire_68, CLK, g1333);
MUX2_X1 g_tmp_wire_69 (g6864, g1333, SE, tmp_wire_69);
DFF_X1 g_g1336 (tmp_wire_69, CLK, g1336);
MUX2_X1 g_tmp_wire_70 (g6865, g1336, SE, tmp_wire_70);
DFF_X1 g_g1339 (tmp_wire_70, CLK, g1339);
MUX2_X1 g_tmp_wire_71 (g7119, g1339, SE, tmp_wire_71);
DFF_X1 g_g1342 (tmp_wire_71, CLK, g1342);
MUX2_X1 g_tmp_wire_72 (g7528, g1342, SE, tmp_wire_72);
DFF_X1 g_g1345 (tmp_wire_72, CLK, g1345);
MUX2_X1 g_tmp_wire_73 (g7529, g1345, SE, tmp_wire_73);
DFF_X1 g_g1348 (tmp_wire_73, CLK, g1348);
MUX2_X1 g_tmp_wire_74 (g7530, g1348, SE, tmp_wire_74);
DFF_X1 g_g1351 (tmp_wire_74, CLK, g1351);
MUX2_X1 g_tmp_wire_75 (g7768, g1351, SE, tmp_wire_75);
DFF_X1 g_g1354 (tmp_wire_75, CLK, g1354);
MUX2_X1 g_tmp_wire_76 (g8675, g1354, SE, tmp_wire_76);
DFF_X1 g_g1357 (tmp_wire_76, CLK, g1357);
MUX2_X1 g_tmp_wire_77 (g8676, g1357, SE, tmp_wire_77);
DFF_X1 g_g1360 (tmp_wire_77, CLK, g1360);
MUX2_X1 g_tmp_wire_78 (g8677, g1360, SE, tmp_wire_78);
DFF_X1 g_g1190 (tmp_wire_78, CLK, g1190);
MUX2_X1 g_tmp_wire_79 (g6373, g1190, SE, tmp_wire_79);
DFF_X1 g_g1191 (tmp_wire_79, CLK, g1191);
MUX2_X1 g_tmp_wire_80 (g1191, g1191, SE, tmp_wire_80);
DFF_X1 g_g1192 (tmp_wire_80, CLK, g1192);
MUX2_X1 g_tmp_wire_81 (g1192, g1192, SE, tmp_wire_81);
DFF_X1 g_g1193 (tmp_wire_81, CLK, g1193);
MUX2_X1 g_tmp_wire_82 (g1193, g1193, SE, tmp_wire_82);
DFF_X1 g_g1194 (tmp_wire_82, CLK, g1194);
MUX2_X1 g_tmp_wire_83 (g6374, g1194, SE, tmp_wire_83);
DFF_X1 g_g1195 (tmp_wire_83, CLK, g1195);
MUX2_X1 g_tmp_wire_84 (g1195, g1195, SE, tmp_wire_84);
DFF_X1 g_g1196 (tmp_wire_84, CLK, g1196);
MUX2_X1 g_tmp_wire_85 (g1196, g1196, SE, tmp_wire_85);
DFF_X1 g_g1197 (tmp_wire_85, CLK, g1197);
MUX2_X1 g_tmp_wire_86 (g1197, g1197, SE, tmp_wire_86);
DFF_X1 g_g1198 (tmp_wire_86, CLK, g1198);
MUX2_X1 g_tmp_wire_87 (g6375, g1198, SE, tmp_wire_87);
DFF_X1 g_g1199 (tmp_wire_87, CLK, g1199);
MUX2_X1 g_tmp_wire_88 (g1199, g1199, SE, tmp_wire_88);
DFF_X1 g_g1200 (tmp_wire_88, CLK, g1200);
MUX2_X1 g_tmp_wire_89 (g1200, g1200, SE, tmp_wire_89);
DFF_X1 g_g1201 (tmp_wire_89, CLK, g1201);
MUX2_X1 g_tmp_wire_90 (g1201, g1201, SE, tmp_wire_90);
DFF_X1 g_g1202 (tmp_wire_90, CLK, g1202);
MUX2_X1 g_tmp_wire_91 (g6376, g1202, SE, tmp_wire_91);
DFF_X1 g_g1203 (tmp_wire_91, CLK, g1203);
MUX2_X1 g_tmp_wire_92 (g1203, g1203, SE, tmp_wire_92);
DFF_X1 g_g1204 (tmp_wire_92, CLK, g1204);
MUX2_X1 g_tmp_wire_93 (g1204, g1204, SE, tmp_wire_93);
DFF_X1 g_g1205 (tmp_wire_93, CLK, g1205);
MUX2_X1 g_tmp_wire_94 (g1205, g1205, SE, tmp_wire_94);
DFF_X1 g_g1206 (tmp_wire_94, CLK, g1206);
MUX2_X1 g_tmp_wire_95 (g2661, g1206, SE, tmp_wire_95);
DFF_X1 g_g1252 (tmp_wire_95, CLK, g1252);
MUX2_X1 g_tmp_wire_96 (g7111, g1252, SE, tmp_wire_96);
DFF_X1 g_g1250 (tmp_wire_96, CLK, g1250);
MUX2_X1 g_tmp_wire_97 (g6860, g1250, SE, tmp_wire_97);
DFF_X1 g_g1251 (tmp_wire_97, CLK, g1251);
MUX2_X1 g_tmp_wire_98 (g6380, g1251, SE, tmp_wire_98);
DFF_X1 g_g1247 (tmp_wire_98, CLK, g1247);
MUX2_X1 g_tmp_wire_99 (g6381, g1247, SE, tmp_wire_99);
DFF_X1 g_g1254 (tmp_wire_99, CLK, g1254);
MUX2_X1 g_tmp_wire_100 (g5739, g1254, SE, tmp_wire_100);
DFF_X1 g_g1266 (tmp_wire_100, CLK, g1266);
MUX2_X1 g_tmp_wire_101 (g6382, g1266, SE, tmp_wire_101);
DFF_X1 g_g1260 (tmp_wire_101, CLK, g1260);
MUX2_X1 g_tmp_wire_102 (g5738, g1260, SE, tmp_wire_102);
DFF_X1 g_g1257 (tmp_wire_102, CLK, g1257);
MUX2_X1 g_tmp_wire_103 (g5737, g1257, SE, tmp_wire_103);
DFF_X1 g_g1263 (tmp_wire_103, CLK, g1263);
MUX2_X1 g_tmp_wire_104 (g4656, g1263, SE, tmp_wire_104);
DFF_X1 g_g1267 (tmp_wire_104, CLK, g1267);
MUX2_X1 g_tmp_wire_105 (g5175, g1267, SE, tmp_wire_105);
DFF_X1 g_g1268 (tmp_wire_105, CLK, g1268);
MUX2_X1 g_tmp_wire_106 (g5740, g1268, SE, tmp_wire_106);
DFF_X1 g_g1269 (tmp_wire_106, CLK, g1269);
MUX2_X1 g_tmp_wire_107 (g5176, g1269, SE, tmp_wire_107);
DFF_X1 g_g1271 (tmp_wire_107, CLK, g1271);
MUX2_X1 g_tmp_wire_108 (g1271, g1271, SE, tmp_wire_108);
DFF_X1 g_g1270 (tmp_wire_108, CLK, g1270);
MUX2_X1 g_tmp_wire_109 (g1270, g1270, SE, tmp_wire_109);
DFF_X1 g_g172 (tmp_wire_109, CLK, g172);
MUX2_X1 g_tmp_wire_110 (g5742, g172, SE, tmp_wire_110);
DFF_X1 g_g1313 (tmp_wire_110, CLK, g1313);
MUX2_X1 g_tmp_wire_111 (g5743, g1313, SE, tmp_wire_111);
DFF_X1 g_g1317 (tmp_wire_111, CLK, g1317);
MUX2_X1 g_tmp_wire_112 (g6861, g1317, SE, tmp_wire_112);
DFF_X1 g_g1318 (tmp_wire_112, CLK, g1318);
MUX2_X1 g_tmp_wire_113 (g7113, g1318, SE, tmp_wire_113);
DFF_X1 g_g1319 (tmp_wire_113, CLK, g1319);
MUX2_X1 g_tmp_wire_114 (g7114, g1319, SE, tmp_wire_114);
DFF_X1 g_g1320 (tmp_wire_114, CLK, g1320);
MUX2_X1 g_tmp_wire_115 (g7115, g1320, SE, tmp_wire_115);
DFF_X1 g_g1321 (tmp_wire_115, CLK, g1321);
MUX2_X1 g_tmp_wire_116 (g7116, g1321, SE, tmp_wire_116);
DFF_X1 g_g1322 (tmp_wire_116, CLK, g1322);
MUX2_X1 g_tmp_wire_117 (g7117, g1322, SE, tmp_wire_117);
DFF_X1 g_g1323 (tmp_wire_117, CLK, g1323);
MUX2_X1 g_tmp_wire_118 (g7118, g1323, SE, tmp_wire_118);
DFF_X1 g_g1324 (tmp_wire_118, CLK, g1324);
MUX2_X1 g_tmp_wire_119 (g7305, g1324, SE, tmp_wire_119);
DFF_X1 g_g1325 (tmp_wire_119, CLK, g1325);
MUX2_X1 g_tmp_wire_120 (g7306, g1325, SE, tmp_wire_120);
DFF_X1 g_g1326 (tmp_wire_120, CLK, g1326);
MUX2_X1 g_tmp_wire_121 (g7307, g1326, SE, tmp_wire_121);
DFF_X1 g_g1327 (tmp_wire_121, CLK, g1327);
MUX2_X1 g_tmp_wire_122 (g7309, g1327, SE, tmp_wire_122);
DFF_X1 g_g1328 (tmp_wire_122, CLK, g1328);
MUX2_X1 g_tmp_wire_123 (g7308, g1328, SE, tmp_wire_123);
DFF_X1 g_g13 (tmp_wire_123, CLK, g13);
MUX2_X1 g_tmp_wire_124 (g2663, g13, SE, tmp_wire_124);
DFF_X1 g_g1329 (tmp_wire_124, CLK, g1329);
MUX2_X1 g_tmp_wire_125 (g6386, g1329, SE, tmp_wire_125);
DFF_X1 g_g20 (tmp_wire_125, CLK, g20);
MUX2_X1 g_tmp_wire_126 (g6866, g20, SE, tmp_wire_126);
DFF_X1 g_g1366 (tmp_wire_126, CLK, g1366);
MUX2_X1 g_tmp_wire_127 (g6878, g1366, SE, tmp_wire_127);
DFF_X1 g_g1364 (tmp_wire_127, CLK, g1364);
MUX2_X1 g_tmp_wire_128 (g6876, g1364, SE, tmp_wire_128);
DFF_X1 g_g1370 (tmp_wire_128, CLK, g1370);
MUX2_X1 g_tmp_wire_129 (g6874, g1370, SE, tmp_wire_129);
DFF_X1 g_g1368 (tmp_wire_129, CLK, g1368);
MUX2_X1 g_tmp_wire_130 (g6872, g1368, SE, tmp_wire_130);
DFF_X1 g_g1374 (tmp_wire_130, CLK, g1374);
MUX2_X1 g_tmp_wire_131 (g6870, g1374, SE, tmp_wire_131);
DFF_X1 g_g1372 (tmp_wire_131, CLK, g1372);
MUX2_X1 g_tmp_wire_132 (g6869, g1372, SE, tmp_wire_132);
DFF_X1 g_g1375 (tmp_wire_132, CLK, g1375);
MUX2_X1 g_tmp_wire_133 (g6867, g1375, SE, tmp_wire_133);
DFF_X1 g_g1365 (tmp_wire_133, CLK, g1365);
MUX2_X1 g_tmp_wire_134 (g6877, g1365, SE, tmp_wire_134);
DFF_X1 g_g1363 (tmp_wire_134, CLK, g1363);
MUX2_X1 g_tmp_wire_135 (g6875, g1363, SE, tmp_wire_135);
DFF_X1 g_g1369 (tmp_wire_135, CLK, g1369);
MUX2_X1 g_tmp_wire_136 (g6873, g1369, SE, tmp_wire_136);
DFF_X1 g_g1367 (tmp_wire_136, CLK, g1367);
MUX2_X1 g_tmp_wire_137 (g6871, g1367, SE, tmp_wire_137);
DFF_X1 g_g1373 (tmp_wire_137, CLK, g1373);
MUX2_X1 g_tmp_wire_138 (g6868, g1373, SE, tmp_wire_138);
DFF_X1 g_g1371 (tmp_wire_138, CLK, g1371);
MUX2_X1 g_tmp_wire_139 (g4658, g1371, SE, tmp_wire_139);
DFF_X1 g_g1389 (tmp_wire_139, CLK, g1389);
MUX2_X1 g_tmp_wire_140 (g6879, g1389, SE, tmp_wire_140);
DFF_X1 g_g1379 (tmp_wire_140, CLK, g1379);
MUX2_X1 g_tmp_wire_141 (g6891, g1379, SE, tmp_wire_141);
DFF_X1 g_g1377 (tmp_wire_141, CLK, g1377);
MUX2_X1 g_tmp_wire_142 (g6889, g1377, SE, tmp_wire_142);
DFF_X1 g_g1383 (tmp_wire_142, CLK, g1383);
MUX2_X1 g_tmp_wire_143 (g6887, g1383, SE, tmp_wire_143);
DFF_X1 g_g1381 (tmp_wire_143, CLK, g1381);
MUX2_X1 g_tmp_wire_144 (g6885, g1381, SE, tmp_wire_144);
DFF_X1 g_g1387 (tmp_wire_144, CLK, g1387);
MUX2_X1 g_tmp_wire_145 (g6883, g1387, SE, tmp_wire_145);
DFF_X1 g_g1385 (tmp_wire_145, CLK, g1385);
MUX2_X1 g_tmp_wire_146 (g6882, g1385, SE, tmp_wire_146);
DFF_X1 g_g1388 (tmp_wire_146, CLK, g1388);
MUX2_X1 g_tmp_wire_147 (g6880, g1388, SE, tmp_wire_147);
DFF_X1 g_g1378 (tmp_wire_147, CLK, g1378);
MUX2_X1 g_tmp_wire_148 (g6890, g1378, SE, tmp_wire_148);
DFF_X1 g_g1376 (tmp_wire_148, CLK, g1376);
MUX2_X1 g_tmp_wire_149 (g6888, g1376, SE, tmp_wire_149);
DFF_X1 g_g1382 (tmp_wire_149, CLK, g1382);
MUX2_X1 g_tmp_wire_150 (g6886, g1382, SE, tmp_wire_150);
DFF_X1 g_g1380 (tmp_wire_150, CLK, g1380);
MUX2_X1 g_tmp_wire_151 (g6884, g1380, SE, tmp_wire_151);
DFF_X1 g_g1386 (tmp_wire_151, CLK, g1386);
MUX2_X1 g_tmp_wire_152 (g6881, g1386, SE, tmp_wire_152);
DFF_X1 g_g1384 (tmp_wire_152, CLK, g1384);
MUX2_X1 g_tmp_wire_153 (g4659, g1384, SE, tmp_wire_153);
DFF_X1 g_g1390 (tmp_wire_153, CLK, g1390);
MUX2_X1 g_tmp_wire_154 (g1390, g1390, SE, tmp_wire_154);
DFF_X1 g_g1391 (tmp_wire_154, CLK, g1391);
MUX2_X1 g_tmp_wire_155 (g6387, g1391, SE, tmp_wire_155);
DFF_X1 g_g1392 (tmp_wire_155, CLK, g1392);
MUX2_X1 g_tmp_wire_156 (g2664, g1392, SE, tmp_wire_156);
DFF_X1 g_g1393 (tmp_wire_156, CLK, g1393);
MUX2_X1 g_tmp_wire_157 (g1393, g1393, SE, tmp_wire_157);
DFF_X1 g_g1395 (tmp_wire_157, CLK, g1395);
MUX2_X1 g_tmp_wire_158 (g6388, g1395, SE, tmp_wire_158);
DFF_X1 g_g1394 (tmp_wire_158, CLK, g1394);
MUX2_X1 g_tmp_wire_159 (g4662, g1394, SE, tmp_wire_159);
DFF_X1 g_g1396 (tmp_wire_159, CLK, g1396);
MUX2_X1 g_tmp_wire_160 (g1396, g1396, SE, tmp_wire_160);
DFF_X1 g_g1398 (tmp_wire_160, CLK, g1398);
MUX2_X1 g_tmp_wire_161 (g6389, g1398, SE, tmp_wire_161);
DFF_X1 g_g1397 (tmp_wire_161, CLK, g1397);
MUX2_X1 g_tmp_wire_162 (g3861, g1397, SE, tmp_wire_162);
DFF_X1 g_g1399 (tmp_wire_162, CLK, g1399);
MUX2_X1 g_tmp_wire_163 (g1399, g1399, SE, tmp_wire_163);
DFF_X1 g_g1401 (tmp_wire_163, CLK, g1401);
MUX2_X1 g_tmp_wire_164 (g6390, g1401, SE, tmp_wire_164);
DFF_X1 g_g1400 (tmp_wire_164, CLK, g1400);
MUX2_X1 g_tmp_wire_165 (g6391, g1400, SE, tmp_wire_165);
DFF_X1 g_g1402 (tmp_wire_165, CLK, g1402);
MUX2_X1 g_tmp_wire_166 (g1402, g1402, SE, tmp_wire_166);
DFF_X1 g_g1403 (tmp_wire_166, CLK, g1403);
MUX2_X1 g_tmp_wire_167 (g1403, g1403, SE, tmp_wire_167);
DFF_X1 g_g1404 (tmp_wire_167, CLK, g1404);
MUX2_X1 g_tmp_wire_168 (g1404, g1404, SE, tmp_wire_168);
DFF_X1 g_g16 (tmp_wire_168, CLK, g16);
MUX2_X1 g_tmp_wire_169 (g6392, g16, SE, tmp_wire_169);
DFF_X1 g_g1189 (tmp_wire_169, CLK, g1189);
MUX2_X1 g_tmp_wire_170 (g5745, g1189, SE, tmp_wire_170);
DFF_X1 g_g1412 (tmp_wire_170, CLK, g1412);
MUX2_X1 g_tmp_wire_171 (g5180, g1412, SE, tmp_wire_171);
DFF_X1 g_g1415 (tmp_wire_171, CLK, g1415);
MUX2_X1 g_tmp_wire_172 (g5178, g1415, SE, tmp_wire_172);
DFF_X1 g_g1409 (tmp_wire_172, CLK, g1409);
MUX2_X1 g_tmp_wire_173 (g4665, g1409, SE, tmp_wire_173);
DFF_X1 g_g1416 (tmp_wire_173, CLK, g1416);
MUX2_X1 g_tmp_wire_174 (g5179, g1416, SE, tmp_wire_174);
DFF_X1 g_g1421 (tmp_wire_174, CLK, g1421);
MUX2_X1 g_tmp_wire_175 (g5744, g1421, SE, tmp_wire_175);
DFF_X1 g_g1405 (tmp_wire_175, CLK, g1405);
MUX2_X1 g_tmp_wire_176 (g5177, g1405, SE, tmp_wire_176);
DFF_X1 g_g1408 (tmp_wire_176, CLK, g1408);
MUX2_X1 g_tmp_wire_177 (g2671, g1408, SE, tmp_wire_177);
DFF_X1 g_g1429 (tmp_wire_177, CLK, g1429);
MUX2_X1 g_tmp_wire_178 (g2672, g1429, SE, tmp_wire_178);
DFF_X1 g_g1428 (tmp_wire_178, CLK, g1428);
MUX2_X1 g_tmp_wire_179 (g2673, g1428, SE, tmp_wire_179);
DFF_X1 g_g1431 (tmp_wire_179, CLK, g1431);
MUX2_X1 g_tmp_wire_180 (g4666, g1431, SE, tmp_wire_180);
DFF_X1 g_g1430 (tmp_wire_180, CLK, g1430);
MUX2_X1 g_tmp_wire_181 (g3862, g1430, SE, tmp_wire_181);
DFF_X1 g_g1424 (tmp_wire_181, CLK, g1424);
MUX2_X1 g_tmp_wire_182 (g6393, g1424, SE, tmp_wire_182);
DFF_X1 g_g1524 (tmp_wire_182, CLK, g1524);
MUX2_X1 g_tmp_wire_183 (g1524, g1524, SE, tmp_wire_183);
DFF_X1 g_g1513 (tmp_wire_183, CLK, g1513);
MUX2_X1 g_tmp_wire_184 (g8226, g1513, SE, tmp_wire_184);
DFF_X1 g_g1486 (tmp_wire_184, CLK, g1486);
MUX2_X1 g_tmp_wire_185 (g7769, g1486, SE, tmp_wire_185);
DFF_X1 g_g1481 (tmp_wire_185, CLK, g1481);
MUX2_X1 g_tmp_wire_186 (g7770, g1481, SE, tmp_wire_186);
DFF_X1 g_g1489 (tmp_wire_186, CLK, g1489);
MUX2_X1 g_tmp_wire_187 (g7771, g1489, SE, tmp_wire_187);
DFF_X1 g_g1494 (tmp_wire_187, CLK, g1494);
MUX2_X1 g_tmp_wire_188 (g7772, g1494, SE, tmp_wire_188);
DFF_X1 g_g1499 (tmp_wire_188, CLK, g1499);
MUX2_X1 g_tmp_wire_189 (g7773, g1499, SE, tmp_wire_189);
DFF_X1 g_g1504 (tmp_wire_189, CLK, g1504);
MUX2_X1 g_tmp_wire_190 (g7774, g1504, SE, tmp_wire_190);
DFF_X1 g_g1509 (tmp_wire_190, CLK, g1509);
MUX2_X1 g_tmp_wire_191 (g7775, g1509, SE, tmp_wire_191);
DFF_X1 g_g1514 (tmp_wire_191, CLK, g1514);
MUX2_X1 g_tmp_wire_192 (g8227, g1514, SE, tmp_wire_192);
DFF_X1 g_g1519 (tmp_wire_192, CLK, g1519);
MUX2_X1 g_tmp_wire_193 (g8678, g1519, SE, tmp_wire_193);
DFF_X1 g_g1462 (tmp_wire_193, CLK, g1462);
MUX2_X1 g_tmp_wire_194 (g8875, g1462, SE, tmp_wire_194);
DFF_X1 g_g1467 (tmp_wire_194, CLK, g1467);
MUX2_X1 g_tmp_wire_195 (g8960, g1467, SE, tmp_wire_195);
DFF_X1 g_g1472 (tmp_wire_195, CLK, g1472);
MUX2_X1 g_tmp_wire_196 (g9036, g1472, SE, tmp_wire_196);
DFF_X1 g_g1477 (tmp_wire_196, CLK, g1477);
MUX2_X1 g_tmp_wire_197 (g8228, g1477, SE, tmp_wire_197);
DFF_X1 g_g727 (tmp_wire_197, CLK, g727);
MUX2_X1 g_tmp_wire_198 (g7781, g727, SE, tmp_wire_198);
DFF_X1 g_g1532 (tmp_wire_198, CLK, g1532);
MUX2_X1 g_tmp_wire_199 (g7776, g1532, SE, tmp_wire_199);
DFF_X1 g_g1528 (tmp_wire_199, CLK, g1528);
MUX2_X1 g_tmp_wire_200 (g7777, g1528, SE, tmp_wire_200);
DFF_X1 g_g1537 (tmp_wire_200, CLK, g1537);
MUX2_X1 g_tmp_wire_201 (g7778, g1537, SE, tmp_wire_201);
DFF_X1 g_g1541 (tmp_wire_201, CLK, g1541);
MUX2_X1 g_tmp_wire_202 (g7779, g1541, SE, tmp_wire_202);
DFF_X1 g_g1545 (tmp_wire_202, CLK, g1545);
MUX2_X1 g_tmp_wire_203 (g7780, g1545, SE, tmp_wire_203);
DFF_X1 g_g1549 (tmp_wire_203, CLK, g1549);
MUX2_X1 g_tmp_wire_204 (g5181, g1549, SE, tmp_wire_204);
DFF_X1 g_g1435 (tmp_wire_204, CLK, g1435);
MUX2_X1 g_tmp_wire_205 (g5182, g1435, SE, tmp_wire_205);
DFF_X1 g_g1439 (tmp_wire_205, CLK, g1439);
MUX2_X1 g_tmp_wire_206 (g5183, g1439, SE, tmp_wire_206);
DFF_X1 g_g1432 (tmp_wire_206, CLK, g1432);
MUX2_X1 g_tmp_wire_207 (g4667, g1432, SE, tmp_wire_207);
DFF_X1 g_g1443 (tmp_wire_207, CLK, g1443);
MUX2_X1 g_tmp_wire_208 (g5184, g1443, SE, tmp_wire_208);
DFF_X1 g_g33 (tmp_wire_208, CLK, g33);
MUX2_X1 g_tmp_wire_209 (g5746, g33, SE, tmp_wire_209);
DFF_X1 g_g38 (tmp_wire_209, CLK, g38);
MUX2_X1 g_tmp_wire_210 (g4669, g38, SE, tmp_wire_210);
DFF_X1 g_g1461 (tmp_wire_210, CLK, g1461);
MUX2_X1 g_tmp_wire_211 (g5185, g1461, SE, tmp_wire_211);
DFF_X1 g_g1444 (tmp_wire_211, CLK, g1444);
MUX2_X1 g_tmp_wire_212 (g5186, g1444, SE, tmp_wire_212);
DFF_X1 g_g1450 (tmp_wire_212, CLK, g1450);
MUX2_X1 g_tmp_wire_213 (g5187, g1450, SE, tmp_wire_213);
DFF_X1 g_g1454 (tmp_wire_213, CLK, g1454);
MUX2_X1 g_tmp_wire_214 (g3863, g1454, SE, tmp_wire_214);
DFF_X1 g_g1459 (tmp_wire_214, CLK, g1459);
MUX2_X1 g_tmp_wire_215 (g4668, g1459, SE, tmp_wire_215);
DFF_X1 g_g1460 (tmp_wire_215, CLK, g1460);
MUX2_X1 g_tmp_wire_216 (g7104, g1460, SE, tmp_wire_216);
DFF_X1 g_g979 (tmp_wire_216, CLK, g979);
MUX2_X1 g_tmp_wire_217 (g8223, g979, SE, tmp_wire_217);
DFF_X1 g_g966 (tmp_wire_217, CLK, g966);
MUX2_X1 g_tmp_wire_218 (g966, g966, SE, tmp_wire_218);
DFF_X1 g_g969 (tmp_wire_218, CLK, g969);
MUX2_X1 g_tmp_wire_219 (g7764, g969, SE, tmp_wire_219);
DFF_X1 g_g963 (tmp_wire_219, CLK, g963);
MUX2_X1 g_tmp_wire_220 (g963, g963, SE, tmp_wire_220);
DFF_X1 g_g970 (tmp_wire_220, CLK, g970);
MUX2_X1 g_tmp_wire_221 (g5171, g970, SE, tmp_wire_221);
DFF_X1 g_g971 (tmp_wire_221, CLK, g971);
MUX2_X1 g_tmp_wire_222 (g2653, g971, SE, tmp_wire_222);
DFF_X1 g_g972 (tmp_wire_222, CLK, g972);
MUX2_X1 g_tmp_wire_223 (g8672, g972, SE, tmp_wire_223);
DFF_X1 g_g973 (tmp_wire_223, CLK, g973);
MUX2_X1 g_tmp_wire_224 (g8864, g973, SE, tmp_wire_224);
DFF_X1 g_g976 (tmp_wire_224, CLK, g976);
MUX2_X1 g_tmp_wire_225 (g9133, g976, SE, tmp_wire_225);
DFF_X1 g_g984 (tmp_wire_225, CLK, g984);
MUX2_X1 g_tmp_wire_226 (g7515, g984, SE, tmp_wire_226);
DFF_X1 g_g985 (tmp_wire_226, CLK, g985);
MUX2_X1 g_tmp_wire_227 (g7516, g985, SE, tmp_wire_227);
DFF_X1 g_g990 (tmp_wire_227, CLK, g990);
MUX2_X1 g_tmp_wire_228 (g7517, g990, SE, tmp_wire_228);
DFF_X1 g_g995 (tmp_wire_228, CLK, g995);
MUX2_X1 g_tmp_wire_229 (g7105, g995, SE, tmp_wire_229);
DFF_X1 g_g1004 (tmp_wire_229, CLK, g1004);
MUX2_X1 g_tmp_wire_230 (g1004, g1004, SE, tmp_wire_230);
DFF_X1 g_g1005 (tmp_wire_230, CLK, g1005);
MUX2_X1 g_tmp_wire_231 (g1005, g1005, SE, tmp_wire_231);
DFF_X1 g_g998 (tmp_wire_231, CLK, g998);
MUX2_X1 g_tmp_wire_232 (g8865, g998, SE, tmp_wire_232);
DFF_X1 g_g999 (tmp_wire_232, CLK, g999);
MUX2_X1 g_tmp_wire_233 (g8867, g999, SE, tmp_wire_233);
DFF_X1 g_g1007 (tmp_wire_233, CLK, g1007);
MUX2_X1 g_tmp_wire_234 (g6851, g1007, SE, tmp_wire_234);
DFF_X1 g_g1012 (tmp_wire_234, CLK, g1012);
MUX2_X1 g_tmp_wire_235 (g1012, g1012, SE, tmp_wire_235);
DFF_X1 g_g1014 (tmp_wire_235, CLK, g1014);
MUX2_X1 g_tmp_wire_236 (g1014, g1014, SE, tmp_wire_236);
DFF_X1 g_g1013 (tmp_wire_236, CLK, g1013);
MUX2_X1 g_tmp_wire_237 (g2654, g1013, SE, tmp_wire_237);
DFF_X1 g_g1029 (tmp_wire_237, CLK, g1029);
MUX2_X1 g_tmp_wire_238 (g8869, g1029, SE, tmp_wire_238);
DFF_X1 g_g1018 (tmp_wire_238, CLK, g1018);
MUX2_X1 g_tmp_wire_239 (g8870, g1018, SE, tmp_wire_239);
DFF_X1 g_g1021 (tmp_wire_239, CLK, g1021);
MUX2_X1 g_tmp_wire_240 (g8871, g1021, SE, tmp_wire_240);
DFF_X1 g_g1025 (tmp_wire_240, CLK, g1025);
MUX2_X1 g_tmp_wire_241 (g9034, g1025, SE, tmp_wire_241);
DFF_X1 g_g1033 (tmp_wire_241, CLK, g1033);
MUX2_X1 g_tmp_wire_242 (g8957, g1033, SE, tmp_wire_242);
DFF_X1 g_g1034 (tmp_wire_242, CLK, g1034);
MUX2_X1 g_tmp_wire_243 (g7518, g1034, SE, tmp_wire_243);
DFF_X1 g_g1030 (tmp_wire_243, CLK, g1030);
MUX2_X1 g_tmp_wire_244 (g6852, g1030, SE, tmp_wire_244);
DFF_X1 g_g1081 (tmp_wire_244, CLK, g1081);
MUX2_X1 g_tmp_wire_245 (g1081, g1081, SE, tmp_wire_245);
DFF_X1 g_g1156 (tmp_wire_245, CLK, g1156);
MUX2_X1 g_tmp_wire_246 (g1156, g1156, SE, tmp_wire_246);
DFF_X1 g_g1157 (tmp_wire_246, CLK, g1157);
MUX2_X1 g_tmp_wire_247 (g1157, g1157, SE, tmp_wire_247);
DFF_X1 g_g1159 (tmp_wire_247, CLK, g1159);
MUX2_X1 g_tmp_wire_248 (g1159, g1159, SE, tmp_wire_248);
DFF_X1 g_g1158 (tmp_wire_248, CLK, g1158);
MUX2_X1 g_tmp_wire_249 (g7106, g1158, SE, tmp_wire_249);
DFF_X1 g_g1084 (tmp_wire_249, CLK, g1084);
MUX2_X1 g_tmp_wire_250 (g1612, g1084, SE, tmp_wire_250);
DFF_X1 g_g1146 (tmp_wire_250, CLK, g1146);
MUX2_X1 g_tmp_wire_251 (g1146, g1146, SE, tmp_wire_251);
DFF_X1 g_g1147 (tmp_wire_251, CLK, g1147);
MUX2_X1 g_tmp_wire_252 (g1147, g1147, SE, tmp_wire_252);
DFF_X1 g_g1148 (tmp_wire_252, CLK, g1148);
MUX2_X1 g_tmp_wire_253 (g6853, g1148, SE, tmp_wire_253);
DFF_X1 g_g1087 (tmp_wire_253, CLK, g1087);
MUX2_X1 g_tmp_wire_254 (g6854, g1087, SE, tmp_wire_254);
DFF_X1 g_g1098 (tmp_wire_254, CLK, g1098);
MUX2_X1 g_tmp_wire_255 (g6855, g1098, SE, tmp_wire_255);
DFF_X1 g_g1102 (tmp_wire_255, CLK, g1102);
MUX2_X1 g_tmp_wire_256 (g7107, g1102, SE, tmp_wire_256);
DFF_X1 g_g1106 (tmp_wire_256, CLK, g1106);
MUX2_X1 g_tmp_wire_257 (g7299, g1106, SE, tmp_wire_257);
DFF_X1 g_g1110 (tmp_wire_257, CLK, g1110);
MUX2_X1 g_tmp_wire_258 (g7521, g1110, SE, tmp_wire_258);
DFF_X1 g_g1114 (tmp_wire_258, CLK, g1114);
MUX2_X1 g_tmp_wire_259 (g7766, g1114, SE, tmp_wire_259);
DFF_X1 g_g1118 (tmp_wire_259, CLK, g1118);
MUX2_X1 g_tmp_wire_260 (g8225, g1118, SE, tmp_wire_260);
DFF_X1 g_g1122 (tmp_wire_260, CLK, g1122);
MUX2_X1 g_tmp_wire_261 (g8674, g1122, SE, tmp_wire_261);
DFF_X1 g_g1126 (tmp_wire_261, CLK, g1126);
MUX2_X1 g_tmp_wire_262 (g8874, g1126, SE, tmp_wire_262);
DFF_X1 g_g1142 (tmp_wire_262, CLK, g1142);
MUX2_X1 g_tmp_wire_263 (g7526, g1142, SE, tmp_wire_263);
DFF_X1 g_g1173 (tmp_wire_263, CLK, g1173);
MUX2_X1 g_tmp_wire_264 (g1173, g1173, SE, tmp_wire_264);
DFF_X1 g_g1170 (tmp_wire_264, CLK, g1170);
MUX2_X1 g_tmp_wire_265 (g1170, g1170, SE, tmp_wire_265);
DFF_X1 g_g1167 (tmp_wire_265, CLK, g1167);
MUX2_X1 g_tmp_wire_266 (g1167, g1167, SE, tmp_wire_266);
DFF_X1 g_g1166 (tmp_wire_266, CLK, g1166);
MUX2_X1 g_tmp_wire_267 (g7767, g1166, SE, tmp_wire_267);
DFF_X1 g_g1077 (tmp_wire_267, CLK, g1077);
MUX2_X1 g_tmp_wire_268 (g6856, g1077, SE, tmp_wire_268);
DFF_X1 g_g1153 (tmp_wire_268, CLK, g1153);
MUX2_X1 g_tmp_wire_269 (g1153, g1153, SE, tmp_wire_269);
DFF_X1 g_g1154 (tmp_wire_269, CLK, g1154);
MUX2_X1 g_tmp_wire_270 (g1154, g1154, SE, tmp_wire_270);
DFF_X1 g_g1155 (tmp_wire_270, CLK, g1155);
MUX2_X1 g_tmp_wire_271 (g1155, g1155, SE, tmp_wire_271);
DFF_X1 g_g1185 (tmp_wire_271, CLK, g1185);
MUX2_X1 g_tmp_wire_272 (g1185, g1185, SE, tmp_wire_272);
DFF_X1 g_g1097 (tmp_wire_272, CLK, g1097);
MUX2_X1 g_tmp_wire_273 (g7520, g1097, SE, tmp_wire_273);
DFF_X1 g_g1092 (tmp_wire_273, CLK, g1092);
MUX2_X1 g_tmp_wire_274 (g7522, g1092, SE, tmp_wire_274);
DFF_X1 g_g1130 (tmp_wire_274, CLK, g1130);
MUX2_X1 g_tmp_wire_275 (g7523, g1130, SE, tmp_wire_275);
DFF_X1 g_g1134 (tmp_wire_275, CLK, g1134);
MUX2_X1 g_tmp_wire_276 (g7524, g1134, SE, tmp_wire_276);
DFF_X1 g_g1138 (tmp_wire_276, CLK, g1138);
MUX2_X1 g_tmp_wire_277 (g7525, g1138, SE, tmp_wire_277);
DFF_X1 g_g1149 (tmp_wire_277, CLK, g1149);
MUX2_X1 g_tmp_wire_278 (g7519, g1149, SE, tmp_wire_278);
DFF_X1 g_g1037 (tmp_wire_278, CLK, g1037);
MUX2_X1 g_tmp_wire_279 (g7765, g1037, SE, tmp_wire_279);
DFF_X1 g_g1041 (tmp_wire_279, CLK, g1041);
MUX2_X1 g_tmp_wire_280 (g8224, g1041, SE, tmp_wire_280);
DFF_X1 g_g1045 (tmp_wire_280, CLK, g1045);
MUX2_X1 g_tmp_wire_281 (g8673, g1045, SE, tmp_wire_281);
DFF_X1 g_g1049 (tmp_wire_281, CLK, g1049);
MUX2_X1 g_tmp_wire_282 (g8873, g1049, SE, tmp_wire_282);
DFF_X1 g_g1053 (tmp_wire_282, CLK, g1053);
MUX2_X1 g_tmp_wire_283 (g8959, g1053, SE, tmp_wire_283);
DFF_X1 g_g1057 (tmp_wire_283, CLK, g1057);
MUX2_X1 g_tmp_wire_284 (g9035, g1057, SE, tmp_wire_284);
DFF_X1 g_g1061 (tmp_wire_284, CLK, g1061);
MUX2_X1 g_tmp_wire_285 (g9117, g1061, SE, tmp_wire_285);
DFF_X1 g_g1065 (tmp_wire_285, CLK, g1065);
MUX2_X1 g_tmp_wire_286 (g9134, g1065, SE, tmp_wire_286);
DFF_X1 g_g1069 (tmp_wire_286, CLK, g1069);
MUX2_X1 g_tmp_wire_287 (g9145, g1069, SE, tmp_wire_287);
DFF_X1 g_g1073 (tmp_wire_287, CLK, g1073);
MUX2_X1 g_tmp_wire_288 (g2655, g1073, SE, tmp_wire_288);
DFF_X1 g_g1163 (tmp_wire_288, CLK, g1163);
MUX2_X1 g_tmp_wire_289 (g1163, g1163, SE, tmp_wire_289);
DFF_X1 g_g1160 (tmp_wire_289, CLK, g1160);
MUX2_X1 g_tmp_wire_290 (g1160, g1160, SE, tmp_wire_290);
DFF_X1 g_g1182 (tmp_wire_290, CLK, g1182);
MUX2_X1 g_tmp_wire_291 (g1182, g1182, SE, tmp_wire_291);
DFF_X1 g_g1186 (tmp_wire_291, CLK, g1186);
MUX2_X1 g_tmp_wire_292 (g1186, g1186, SE, tmp_wire_292);
DFF_X1 g_g1179 (tmp_wire_292, CLK, g1179);
MUX2_X1 g_tmp_wire_293 (g5172, g1179, SE, tmp_wire_293);
DFF_X1 g_g1176 (tmp_wire_293, CLK, g1176);
MUX2_X1 g_tmp_wire_294 (g6774, g1176, SE, tmp_wire_294);
DFF_X1 g_g68 (tmp_wire_294, CLK, g68);
MUX2_X1 g_tmp_wire_295 (g6775, g68, SE, tmp_wire_295);
DFF_X1 g_g71 (tmp_wire_295, CLK, g71);
MUX2_X1 g_tmp_wire_296 (g6776, g71, SE, tmp_wire_296);
DFF_X1 g_g74 (tmp_wire_296, CLK, g74);
MUX2_X1 g_tmp_wire_297 (g6777, g74, SE, tmp_wire_297);
DFF_X1 g_g77 (tmp_wire_297, CLK, g77);
MUX2_X1 g_tmp_wire_298 (g6778, g77, SE, tmp_wire_298);
DFF_X1 g_g80 (tmp_wire_298, CLK, g80);
MUX2_X1 g_tmp_wire_299 (g6779, g80, SE, tmp_wire_299);
DFF_X1 g_g83 (tmp_wire_299, CLK, g83);
MUX2_X1 g_tmp_wire_300 (g6780, g83, SE, tmp_wire_300);
DFF_X1 g_g86 (tmp_wire_300, CLK, g86);
MUX2_X1 g_tmp_wire_301 (g6781, g86, SE, tmp_wire_301);
DFF_X1 g_g52 (tmp_wire_301, CLK, g52);
MUX2_X1 g_tmp_wire_302 (g7733, g52, SE, tmp_wire_302);
DFF_X1 g_g55 (tmp_wire_302, CLK, g55);
MUX2_X1 g_tmp_wire_303 (g7509, g55, SE, tmp_wire_303);
DFF_X1 g_g62 (tmp_wire_303, CLK, g62);
MUX2_X1 g_tmp_wire_304 (g7734, g62, SE, tmp_wire_304);
DFF_X1 g_g58 (tmp_wire_304, CLK, g58);
MUX2_X1 g_tmp_wire_305 (g4598, g58, SE, tmp_wire_305);
DFF_X1 g_g65 (tmp_wire_305, CLK, g65);
MUX2_X1 g_tmp_wire_306 (g3832, g65, SE, tmp_wire_306);
DFF_X1 g_g199 (tmp_wire_306, CLK, g199);
MUX2_X1 g_tmp_wire_307 (g199, g199, SE, tmp_wire_307);
DFF_X1 g_g200 (tmp_wire_307, CLK, g200);
MUX2_X1 g_tmp_wire_308 (g200, g200, SE, tmp_wire_308);
DFF_X1 g_g201 (tmp_wire_308, CLK, g201);
MUX2_X1 g_tmp_wire_309 (g201, g201, SE, tmp_wire_309);
DFF_X1 g_g190 (tmp_wire_309, CLK, g190);
MUX2_X1 g_tmp_wire_310 (g3831, g190, SE, tmp_wire_310);
DFF_X1 g_g195 (tmp_wire_310, CLK, g195);
MUX2_X1 g_tmp_wire_311 (g5731, g195, SE, tmp_wire_311);
DFF_X1 g_g196 (tmp_wire_311, CLK, g196);
MUX2_X1 g_tmp_wire_312 (g5159, g196, SE, tmp_wire_312);
DFF_X1 g_g179 (tmp_wire_312, CLK, g179);
MUX2_X1 g_tmp_wire_313 (g3830, g179, SE, tmp_wire_313);
DFF_X1 g_g186 (tmp_wire_313, CLK, g186);
MUX2_X1 g_tmp_wire_314 (g5730, g186, SE, tmp_wire_314);
DFF_X1 g_g187 (tmp_wire_314, CLK, g187);
MUX2_X1 g_tmp_wire_315 (g5158, g187, SE, tmp_wire_315);
DFF_X1 g_g180 (tmp_wire_315, CLK, g180);
MUX2_X1 g_tmp_wire_316 (g3835, g180, SE, tmp_wire_316);
DFF_X1 g_g205 (tmp_wire_316, CLK, g205);
MUX2_X1 g_tmp_wire_317 (g5732, g205, SE, tmp_wire_317);
DFF_X1 g_g202 (tmp_wire_317, CLK, g202);
MUX2_X1 g_tmp_wire_318 (g5160, g202, SE, tmp_wire_318);
DFF_X1 g_g181 (tmp_wire_318, CLK, g181);
MUX2_X1 g_tmp_wire_319 (g3834, g181, SE, tmp_wire_319);
DFF_X1 g_g210 (tmp_wire_319, CLK, g210);
MUX2_X1 g_tmp_wire_320 (g5733, g210, SE, tmp_wire_320);
DFF_X1 g_g207 (tmp_wire_320, CLK, g207);
MUX2_X1 g_tmp_wire_321 (g5161, g207, SE, tmp_wire_321);
DFF_X1 g_g182 (tmp_wire_321, CLK, g182);
MUX2_X1 g_tmp_wire_322 (g7735, g182, SE, tmp_wire_322);
DFF_X1 g_g146 (tmp_wire_322, CLK, g146);
MUX2_X1 g_tmp_wire_323 (g7736, g146, SE, tmp_wire_323);
DFF_X1 g_g173 (tmp_wire_323, CLK, g173);
MUX2_X1 g_tmp_wire_324 (g7738, g173, SE, tmp_wire_324);
DFF_X1 g_g150 (tmp_wire_324, CLK, g150);
MUX2_X1 g_tmp_wire_325 (g7737, g150, SE, tmp_wire_325);
DFF_X1 g_g174 (tmp_wire_325, CLK, g174);
MUX2_X1 g_tmp_wire_326 (g7739, g174, SE, tmp_wire_326);
DFF_X1 g_g154 (tmp_wire_326, CLK, g154);
MUX2_X1 g_tmp_wire_327 (g7740, g154, SE, tmp_wire_327);
DFF_X1 g_g158 (tmp_wire_327, CLK, g158);
MUX2_X1 g_tmp_wire_328 (g7741, g158, SE, tmp_wire_328);
DFF_X1 g_g162 (tmp_wire_328, CLK, g162);
MUX2_X1 g_tmp_wire_329 (g7742, g162, SE, tmp_wire_329);
DFF_X1 g_g168 (tmp_wire_329, CLK, g168);
MUX2_X1 g_tmp_wire_330 (g6309, g168, SE, tmp_wire_330);
DFF_X1 g_g183 (tmp_wire_330, CLK, g183);
MUX2_X1 g_tmp_wire_331 (g6310, g183, SE, tmp_wire_331);
DFF_X1 g_g184 (tmp_wire_331, CLK, g184);
MUX2_X1 g_tmp_wire_332 (g4599, g184, SE, tmp_wire_332);
DFF_X1 g_g185 (tmp_wire_332, CLK, g185);
MUX2_X1 g_tmp_wire_333 (g6794, g185, SE, tmp_wire_333);
DFF_X1 g_g92 (tmp_wire_333, CLK, g92);
MUX2_X1 g_tmp_wire_334 (g92, g92, SE, tmp_wire_334);
DFF_X1 g_g89 (tmp_wire_334, CLK, g89);
MUX2_X1 g_tmp_wire_335 (g5145, g89, SE, tmp_wire_335);
DFF_X1 g_g93 (tmp_wire_335, CLK, g93);
MUX2_X1 g_tmp_wire_336 (g6782, g93, SE, tmp_wire_336);
DFF_X1 g_g94 (tmp_wire_336, CLK, g94);
MUX2_X1 g_tmp_wire_337 (g94, g94, SE, tmp_wire_337);
DFF_X1 g_g95 (tmp_wire_337, CLK, g95);
MUX2_X1 g_tmp_wire_338 (g5146, g95, SE, tmp_wire_338);
DFF_X1 g_g98 (tmp_wire_338, CLK, g98);
MUX2_X1 g_tmp_wire_339 (g6783, g98, SE, tmp_wire_339);
DFF_X1 g_g99 (tmp_wire_339, CLK, g99);
MUX2_X1 g_tmp_wire_340 (g99, g99, SE, tmp_wire_340);
DFF_X1 g_g100 (tmp_wire_340, CLK, g100);
MUX2_X1 g_tmp_wire_341 (g5157, g100, SE, tmp_wire_341);
DFF_X1 g_g103 (tmp_wire_341, CLK, g103);
MUX2_X1 g_tmp_wire_342 (g6784, g103, SE, tmp_wire_342);
DFF_X1 g_g104 (tmp_wire_342, CLK, g104);
MUX2_X1 g_tmp_wire_343 (g104, g104, SE, tmp_wire_343);
DFF_X1 g_g105 (tmp_wire_343, CLK, g105);
MUX2_X1 g_tmp_wire_344 (g5147, g105, SE, tmp_wire_344);
DFF_X1 g_g108 (tmp_wire_344, CLK, g108);
MUX2_X1 g_tmp_wire_345 (g6785, g108, SE, tmp_wire_345);
DFF_X1 g_g109 (tmp_wire_345, CLK, g109);
MUX2_X1 g_tmp_wire_346 (g109, g109, SE, tmp_wire_346);
DFF_X1 g_g110 (tmp_wire_346, CLK, g110);
MUX2_X1 g_tmp_wire_347 (g5148, g110, SE, tmp_wire_347);
DFF_X1 g_g113 (tmp_wire_347, CLK, g113);
MUX2_X1 g_tmp_wire_348 (g6786, g113, SE, tmp_wire_348);
DFF_X1 g_g114 (tmp_wire_348, CLK, g114);
MUX2_X1 g_tmp_wire_349 (g5153, g114, SE, tmp_wire_349);
DFF_X1 g_g117 (tmp_wire_349, CLK, g117);
MUX2_X1 g_tmp_wire_350 (g6787, g117, SE, tmp_wire_350);
DFF_X1 g_g118 (tmp_wire_350, CLK, g118);
MUX2_X1 g_tmp_wire_351 (g5154, g118, SE, tmp_wire_351);
DFF_X1 g_g121 (tmp_wire_351, CLK, g121);
MUX2_X1 g_tmp_wire_352 (g6788, g121, SE, tmp_wire_352);
DFF_X1 g_g122 (tmp_wire_352, CLK, g122);
MUX2_X1 g_tmp_wire_353 (g5155, g122, SE, tmp_wire_353);
DFF_X1 g_g125 (tmp_wire_353, CLK, g125);
MUX2_X1 g_tmp_wire_354 (g6789, g125, SE, tmp_wire_354);
DFF_X1 g_g126 (tmp_wire_354, CLK, g126);
MUX2_X1 g_tmp_wire_355 (g5156, g126, SE, tmp_wire_355);
DFF_X1 g_g129 (tmp_wire_355, CLK, g129);
MUX2_X1 g_tmp_wire_356 (g6790, g129, SE, tmp_wire_356);
DFF_X1 g_g130 (tmp_wire_356, CLK, g130);
MUX2_X1 g_tmp_wire_357 (g5149, g130, SE, tmp_wire_357);
DFF_X1 g_g133 (tmp_wire_357, CLK, g133);
MUX2_X1 g_tmp_wire_358 (g6791, g133, SE, tmp_wire_358);
DFF_X1 g_g134 (tmp_wire_358, CLK, g134);
MUX2_X1 g_tmp_wire_359 (g5150, g134, SE, tmp_wire_359);
DFF_X1 g_g137 (tmp_wire_359, CLK, g137);
MUX2_X1 g_tmp_wire_360 (g6792, g137, SE, tmp_wire_360);
DFF_X1 g_g138 (tmp_wire_360, CLK, g138);
MUX2_X1 g_tmp_wire_361 (g5151, g138, SE, tmp_wire_361);
DFF_X1 g_g141 (tmp_wire_361, CLK, g141);
MUX2_X1 g_tmp_wire_362 (g6793, g141, SE, tmp_wire_362);
DFF_X1 g_g142 (tmp_wire_362, CLK, g142);
MUX2_X1 g_tmp_wire_363 (g5152, g142, SE, tmp_wire_363);
DFF_X1 g_g145 (tmp_wire_363, CLK, g145);
MUX2_X1 g_tmp_wire_364 (g3836, g145, SE, tmp_wire_364);
DFF_X1 g_g287 (tmp_wire_364, CLK, g287);
MUX2_X1 g_tmp_wire_365 (g287, g287, SE, tmp_wire_365);
DFF_X1 g_g290 (tmp_wire_365, CLK, g290);
MUX2_X1 g_tmp_wire_366 (g9087, g290, SE, tmp_wire_366);
DFF_X1 g_g255 (tmp_wire_366, CLK, g255);
MUX2_X1 g_tmp_wire_367 (g9088, g255, SE, tmp_wire_367);
DFF_X1 g_g258 (tmp_wire_367, CLK, g258);
MUX2_X1 g_tmp_wire_368 (g9089, g258, SE, tmp_wire_368);
DFF_X1 g_g261 (tmp_wire_368, CLK, g261);
MUX2_X1 g_tmp_wire_369 (g9090, g261, SE, tmp_wire_369);
DFF_X1 g_g264 (tmp_wire_369, CLK, g264);
MUX2_X1 g_tmp_wire_370 (g9091, g264, SE, tmp_wire_370);
DFF_X1 g_g267 (tmp_wire_370, CLK, g267);
MUX2_X1 g_tmp_wire_371 (g9092, g267, SE, tmp_wire_371);
DFF_X1 g_g270 (tmp_wire_371, CLK, g270);
MUX2_X1 g_tmp_wire_372 (g9085, g270, SE, tmp_wire_372);
DFF_X1 g_g281 (tmp_wire_372, CLK, g281);
MUX2_X1 g_tmp_wire_373 (g9086, g281, SE, tmp_wire_373);
DFF_X1 g_g284 (tmp_wire_373, CLK, g284);
MUX2_X1 g_tmp_wire_374 (g4600, g284, SE, tmp_wire_374);
DFF_X1 g_g211 (tmp_wire_374, CLK, g211);
MUX2_X1 g_tmp_wire_375 (g6311, g211, SE, tmp_wire_375);
DFF_X1 g_g216 (tmp_wire_375, CLK, g216);
MUX2_X1 g_tmp_wire_376 (g4601, g216, SE, tmp_wire_376);
DFF_X1 g_g212 (tmp_wire_376, CLK, g212);
MUX2_X1 g_tmp_wire_377 (g6312, g212, SE, tmp_wire_377);
DFF_X1 g_g219 (tmp_wire_377, CLK, g219);
MUX2_X1 g_tmp_wire_378 (g4602, g219, SE, tmp_wire_378);
DFF_X1 g_g213 (tmp_wire_378, CLK, g213);
MUX2_X1 g_tmp_wire_379 (g6313, g213, SE, tmp_wire_379);
DFF_X1 g_g222 (tmp_wire_379, CLK, g222);
MUX2_X1 g_tmp_wire_380 (g4603, g222, SE, tmp_wire_380);
DFF_X1 g_g214 (tmp_wire_380, CLK, g214);
MUX2_X1 g_tmp_wire_381 (g6314, g214, SE, tmp_wire_381);
DFF_X1 g_g225 (tmp_wire_381, CLK, g225);
MUX2_X1 g_tmp_wire_382 (g4604, g225, SE, tmp_wire_382);
DFF_X1 g_g215 (tmp_wire_382, CLK, g215);
MUX2_X1 g_tmp_wire_383 (g6315, g215, SE, tmp_wire_383);
DFF_X1 g_g228 (tmp_wire_383, CLK, g228);
MUX2_X1 g_tmp_wire_384 (g4605, g228, SE, tmp_wire_384);
DFF_X1 g_g231 (tmp_wire_384, CLK, g231);
MUX2_X1 g_tmp_wire_385 (g6316, g231, SE, tmp_wire_385);
DFF_X1 g_g237 (tmp_wire_385, CLK, g237);
MUX2_X1 g_tmp_wire_386 (g4606, g237, SE, tmp_wire_386);
DFF_X1 g_g232 (tmp_wire_386, CLK, g232);
MUX2_X1 g_tmp_wire_387 (g6317, g232, SE, tmp_wire_387);
DFF_X1 g_g240 (tmp_wire_387, CLK, g240);
MUX2_X1 g_tmp_wire_388 (g4607, g240, SE, tmp_wire_388);
DFF_X1 g_g233 (tmp_wire_388, CLK, g233);
MUX2_X1 g_tmp_wire_389 (g6318, g233, SE, tmp_wire_389);
DFF_X1 g_g243 (tmp_wire_389, CLK, g243);
MUX2_X1 g_tmp_wire_390 (g4608, g243, SE, tmp_wire_390);
DFF_X1 g_g234 (tmp_wire_390, CLK, g234);
MUX2_X1 g_tmp_wire_391 (g6319, g234, SE, tmp_wire_391);
DFF_X1 g_g246 (tmp_wire_391, CLK, g246);
MUX2_X1 g_tmp_wire_392 (g4609, g246, SE, tmp_wire_392);
DFF_X1 g_g235 (tmp_wire_392, CLK, g235);
MUX2_X1 g_tmp_wire_393 (g6320, g235, SE, tmp_wire_393);
DFF_X1 g_g249 (tmp_wire_393, CLK, g249);
MUX2_X1 g_tmp_wire_394 (g4610, g249, SE, tmp_wire_394);
DFF_X1 g_g236 (tmp_wire_394, CLK, g236);
MUX2_X1 g_tmp_wire_395 (g6321, g236, SE, tmp_wire_395);
DFF_X1 g_g252 (tmp_wire_395, CLK, g252);
MUX2_X1 g_tmp_wire_396 (g4611, g252, SE, tmp_wire_396);
DFF_X1 g_g273 (tmp_wire_396, CLK, g273);
MUX2_X1 g_tmp_wire_397 (g6322, g273, SE, tmp_wire_397);
DFF_X1 g_g275 (tmp_wire_397, CLK, g275);
MUX2_X1 g_tmp_wire_398 (g4612, g275, SE, tmp_wire_398);
DFF_X1 g_g274 (tmp_wire_398, CLK, g274);
MUX2_X1 g_tmp_wire_399 (g6323, g274, SE, tmp_wire_399);
DFF_X1 g_g278 (tmp_wire_399, CLK, g278);
MUX2_X1 g_tmp_wire_400 (g3838, g278, SE, tmp_wire_400);
DFF_X1 g_g368 (tmp_wire_400, CLK, g368);
MUX2_X1 g_tmp_wire_401 (g368, g368, SE, tmp_wire_401);
DFF_X1 g_g371 (tmp_wire_401, CLK, g371);
MUX2_X1 g_tmp_wire_402 (g9095, g371, SE, tmp_wire_402);
DFF_X1 g_g336 (tmp_wire_402, CLK, g336);
MUX2_X1 g_tmp_wire_403 (g9096, g336, SE, tmp_wire_403);
DFF_X1 g_g339 (tmp_wire_403, CLK, g339);
MUX2_X1 g_tmp_wire_404 (g9097, g339, SE, tmp_wire_404);
DFF_X1 g_g342 (tmp_wire_404, CLK, g342);
MUX2_X1 g_tmp_wire_405 (g9098, g342, SE, tmp_wire_405);
DFF_X1 g_g345 (tmp_wire_405, CLK, g345);
MUX2_X1 g_tmp_wire_406 (g9099, g345, SE, tmp_wire_406);
DFF_X1 g_g348 (tmp_wire_406, CLK, g348);
MUX2_X1 g_tmp_wire_407 (g9100, g348, SE, tmp_wire_407);
DFF_X1 g_g351 (tmp_wire_407, CLK, g351);
MUX2_X1 g_tmp_wire_408 (g9093, g351, SE, tmp_wire_408);
DFF_X1 g_g362 (tmp_wire_408, CLK, g362);
MUX2_X1 g_tmp_wire_409 (g9094, g362, SE, tmp_wire_409);
DFF_X1 g_g365 (tmp_wire_409, CLK, g365);
MUX2_X1 g_tmp_wire_410 (g4613, g365, SE, tmp_wire_410);
DFF_X1 g_g292 (tmp_wire_410, CLK, g292);
MUX2_X1 g_tmp_wire_411 (g6324, g292, SE, tmp_wire_411);
DFF_X1 g_g297 (tmp_wire_411, CLK, g297);
MUX2_X1 g_tmp_wire_412 (g4614, g297, SE, tmp_wire_412);
DFF_X1 g_g293 (tmp_wire_412, CLK, g293);
MUX2_X1 g_tmp_wire_413 (g6325, g293, SE, tmp_wire_413);
DFF_X1 g_g300 (tmp_wire_413, CLK, g300);
MUX2_X1 g_tmp_wire_414 (g4615, g300, SE, tmp_wire_414);
DFF_X1 g_g294 (tmp_wire_414, CLK, g294);
MUX2_X1 g_tmp_wire_415 (g6326, g294, SE, tmp_wire_415);
DFF_X1 g_g303 (tmp_wire_415, CLK, g303);
MUX2_X1 g_tmp_wire_416 (g4616, g303, SE, tmp_wire_416);
DFF_X1 g_g295 (tmp_wire_416, CLK, g295);
MUX2_X1 g_tmp_wire_417 (g6327, g295, SE, tmp_wire_417);
DFF_X1 g_g306 (tmp_wire_417, CLK, g306);
MUX2_X1 g_tmp_wire_418 (g4617, g306, SE, tmp_wire_418);
DFF_X1 g_g296 (tmp_wire_418, CLK, g296);
MUX2_X1 g_tmp_wire_419 (g6328, g296, SE, tmp_wire_419);
DFF_X1 g_g309 (tmp_wire_419, CLK, g309);
MUX2_X1 g_tmp_wire_420 (g4618, g309, SE, tmp_wire_420);
DFF_X1 g_g312 (tmp_wire_420, CLK, g312);
MUX2_X1 g_tmp_wire_421 (g6329, g312, SE, tmp_wire_421);
DFF_X1 g_g318 (tmp_wire_421, CLK, g318);
MUX2_X1 g_tmp_wire_422 (g4619, g318, SE, tmp_wire_422);
DFF_X1 g_g313 (tmp_wire_422, CLK, g313);
MUX2_X1 g_tmp_wire_423 (g6330, g313, SE, tmp_wire_423);
DFF_X1 g_g321 (tmp_wire_423, CLK, g321);
MUX2_X1 g_tmp_wire_424 (g4620, g321, SE, tmp_wire_424);
DFF_X1 g_g314 (tmp_wire_424, CLK, g314);
MUX2_X1 g_tmp_wire_425 (g6331, g314, SE, tmp_wire_425);
DFF_X1 g_g324 (tmp_wire_425, CLK, g324);
MUX2_X1 g_tmp_wire_426 (g4621, g324, SE, tmp_wire_426);
DFF_X1 g_g315 (tmp_wire_426, CLK, g315);
MUX2_X1 g_tmp_wire_427 (g6332, g315, SE, tmp_wire_427);
DFF_X1 g_g327 (tmp_wire_427, CLK, g327);
MUX2_X1 g_tmp_wire_428 (g4622, g327, SE, tmp_wire_428);
DFF_X1 g_g316 (tmp_wire_428, CLK, g316);
MUX2_X1 g_tmp_wire_429 (g6333, g316, SE, tmp_wire_429);
DFF_X1 g_g330 (tmp_wire_429, CLK, g330);
MUX2_X1 g_tmp_wire_430 (g4623, g330, SE, tmp_wire_430);
DFF_X1 g_g317 (tmp_wire_430, CLK, g317);
MUX2_X1 g_tmp_wire_431 (g6334, g317, SE, tmp_wire_431);
DFF_X1 g_g333 (tmp_wire_431, CLK, g333);
MUX2_X1 g_tmp_wire_432 (g4624, g333, SE, tmp_wire_432);
DFF_X1 g_g354 (tmp_wire_432, CLK, g354);
MUX2_X1 g_tmp_wire_433 (g6335, g354, SE, tmp_wire_433);
DFF_X1 g_g356 (tmp_wire_433, CLK, g356);
MUX2_X1 g_tmp_wire_434 (g4625, g356, SE, tmp_wire_434);
DFF_X1 g_g355 (tmp_wire_434, CLK, g355);
MUX2_X1 g_tmp_wire_435 (g6336, g355, SE, tmp_wire_435);
DFF_X1 g_g359 (tmp_wire_435, CLK, g359);
MUX2_X1 g_tmp_wire_436 (g3840, g359, SE, tmp_wire_436);
DFF_X1 g_g449 (tmp_wire_436, CLK, g449);
MUX2_X1 g_tmp_wire_437 (g449, g449, SE, tmp_wire_437);
DFF_X1 g_g452 (tmp_wire_437, CLK, g452);
MUX2_X1 g_tmp_wire_438 (g9103, g452, SE, tmp_wire_438);
DFF_X1 g_g417 (tmp_wire_438, CLK, g417);
MUX2_X1 g_tmp_wire_439 (g9104, g417, SE, tmp_wire_439);
DFF_X1 g_g420 (tmp_wire_439, CLK, g420);
MUX2_X1 g_tmp_wire_440 (g9105, g420, SE, tmp_wire_440);
DFF_X1 g_g423 (tmp_wire_440, CLK, g423);
MUX2_X1 g_tmp_wire_441 (g9106, g423, SE, tmp_wire_441);
DFF_X1 g_g426 (tmp_wire_441, CLK, g426);
MUX2_X1 g_tmp_wire_442 (g9107, g426, SE, tmp_wire_442);
DFF_X1 g_g429 (tmp_wire_442, CLK, g429);
MUX2_X1 g_tmp_wire_443 (g9108, g429, SE, tmp_wire_443);
DFF_X1 g_g432 (tmp_wire_443, CLK, g432);
MUX2_X1 g_tmp_wire_444 (g9101, g432, SE, tmp_wire_444);
DFF_X1 g_g443 (tmp_wire_444, CLK, g443);
MUX2_X1 g_tmp_wire_445 (g9102, g443, SE, tmp_wire_445);
DFF_X1 g_g446 (tmp_wire_445, CLK, g446);
MUX2_X1 g_tmp_wire_446 (g4626, g446, SE, tmp_wire_446);
DFF_X1 g_g373 (tmp_wire_446, CLK, g373);
MUX2_X1 g_tmp_wire_447 (g6337, g373, SE, tmp_wire_447);
DFF_X1 g_g378 (tmp_wire_447, CLK, g378);
MUX2_X1 g_tmp_wire_448 (g4627, g378, SE, tmp_wire_448);
DFF_X1 g_g374 (tmp_wire_448, CLK, g374);
MUX2_X1 g_tmp_wire_449 (g6338, g374, SE, tmp_wire_449);
DFF_X1 g_g381 (tmp_wire_449, CLK, g381);
MUX2_X1 g_tmp_wire_450 (g4628, g381, SE, tmp_wire_450);
DFF_X1 g_g375 (tmp_wire_450, CLK, g375);
MUX2_X1 g_tmp_wire_451 (g6339, g375, SE, tmp_wire_451);
DFF_X1 g_g384 (tmp_wire_451, CLK, g384);
MUX2_X1 g_tmp_wire_452 (g4629, g384, SE, tmp_wire_452);
DFF_X1 g_g376 (tmp_wire_452, CLK, g376);
MUX2_X1 g_tmp_wire_453 (g6340, g376, SE, tmp_wire_453);
DFF_X1 g_g387 (tmp_wire_453, CLK, g387);
MUX2_X1 g_tmp_wire_454 (g4630, g387, SE, tmp_wire_454);
DFF_X1 g_g377 (tmp_wire_454, CLK, g377);
MUX2_X1 g_tmp_wire_455 (g6341, g377, SE, tmp_wire_455);
DFF_X1 g_g390 (tmp_wire_455, CLK, g390);
MUX2_X1 g_tmp_wire_456 (g4631, g390, SE, tmp_wire_456);
DFF_X1 g_g393 (tmp_wire_456, CLK, g393);
MUX2_X1 g_tmp_wire_457 (g6342, g393, SE, tmp_wire_457);
DFF_X1 g_g399 (tmp_wire_457, CLK, g399);
MUX2_X1 g_tmp_wire_458 (g4632, g399, SE, tmp_wire_458);
DFF_X1 g_g394 (tmp_wire_458, CLK, g394);
MUX2_X1 g_tmp_wire_459 (g6343, g394, SE, tmp_wire_459);
DFF_X1 g_g402 (tmp_wire_459, CLK, g402);
MUX2_X1 g_tmp_wire_460 (g4633, g402, SE, tmp_wire_460);
DFF_X1 g_g395 (tmp_wire_460, CLK, g395);
MUX2_X1 g_tmp_wire_461 (g6344, g395, SE, tmp_wire_461);
DFF_X1 g_g405 (tmp_wire_461, CLK, g405);
MUX2_X1 g_tmp_wire_462 (g4634, g405, SE, tmp_wire_462);
DFF_X1 g_g396 (tmp_wire_462, CLK, g396);
MUX2_X1 g_tmp_wire_463 (g6345, g396, SE, tmp_wire_463);
DFF_X1 g_g408 (tmp_wire_463, CLK, g408);
MUX2_X1 g_tmp_wire_464 (g4635, g408, SE, tmp_wire_464);
DFF_X1 g_g397 (tmp_wire_464, CLK, g397);
MUX2_X1 g_tmp_wire_465 (g6346, g397, SE, tmp_wire_465);
DFF_X1 g_g411 (tmp_wire_465, CLK, g411);
MUX2_X1 g_tmp_wire_466 (g4636, g411, SE, tmp_wire_466);
DFF_X1 g_g398 (tmp_wire_466, CLK, g398);
MUX2_X1 g_tmp_wire_467 (g6347, g398, SE, tmp_wire_467);
DFF_X1 g_g414 (tmp_wire_467, CLK, g414);
MUX2_X1 g_tmp_wire_468 (g4637, g414, SE, tmp_wire_468);
DFF_X1 g_g435 (tmp_wire_468, CLK, g435);
MUX2_X1 g_tmp_wire_469 (g6348, g435, SE, tmp_wire_469);
DFF_X1 g_g437 (tmp_wire_469, CLK, g437);
MUX2_X1 g_tmp_wire_470 (g4638, g437, SE, tmp_wire_470);
DFF_X1 g_g436 (tmp_wire_470, CLK, g436);
MUX2_X1 g_tmp_wire_471 (g6349, g436, SE, tmp_wire_471);
DFF_X1 g_g440 (tmp_wire_471, CLK, g440);
MUX2_X1 g_tmp_wire_472 (g3842, g440, SE, tmp_wire_472);
DFF_X1 g_g530 (tmp_wire_472, CLK, g530);
MUX2_X1 g_tmp_wire_473 (g530, g530, SE, tmp_wire_473);
DFF_X1 g_g533 (tmp_wire_473, CLK, g533);
MUX2_X1 g_tmp_wire_474 (g9111, g533, SE, tmp_wire_474);
DFF_X1 g_g498 (tmp_wire_474, CLK, g498);
MUX2_X1 g_tmp_wire_475 (g9112, g498, SE, tmp_wire_475);
DFF_X1 g_g501 (tmp_wire_475, CLK, g501);
MUX2_X1 g_tmp_wire_476 (g9113, g501, SE, tmp_wire_476);
DFF_X1 g_g504 (tmp_wire_476, CLK, g504);
MUX2_X1 g_tmp_wire_477 (g9114, g504, SE, tmp_wire_477);
DFF_X1 g_g507 (tmp_wire_477, CLK, g507);
MUX2_X1 g_tmp_wire_478 (g9115, g507, SE, tmp_wire_478);
DFF_X1 g_g510 (tmp_wire_478, CLK, g510);
MUX2_X1 g_tmp_wire_479 (g9116, g510, SE, tmp_wire_479);
DFF_X1 g_g513 (tmp_wire_479, CLK, g513);
MUX2_X1 g_tmp_wire_480 (g9109, g513, SE, tmp_wire_480);
DFF_X1 g_g524 (tmp_wire_480, CLK, g524);
MUX2_X1 g_tmp_wire_481 (g9110, g524, SE, tmp_wire_481);
DFF_X1 g_g527 (tmp_wire_481, CLK, g527);
MUX2_X1 g_tmp_wire_482 (g4639, g527, SE, tmp_wire_482);
DFF_X1 g_g454 (tmp_wire_482, CLK, g454);
MUX2_X1 g_tmp_wire_483 (g6350, g454, SE, tmp_wire_483);
DFF_X1 g_g459 (tmp_wire_483, CLK, g459);
MUX2_X1 g_tmp_wire_484 (g4640, g459, SE, tmp_wire_484);
DFF_X1 g_g455 (tmp_wire_484, CLK, g455);
MUX2_X1 g_tmp_wire_485 (g6351, g455, SE, tmp_wire_485);
DFF_X1 g_g462 (tmp_wire_485, CLK, g462);
MUX2_X1 g_tmp_wire_486 (g4641, g462, SE, tmp_wire_486);
DFF_X1 g_g456 (tmp_wire_486, CLK, g456);
MUX2_X1 g_tmp_wire_487 (g6352, g456, SE, tmp_wire_487);
DFF_X1 g_g465 (tmp_wire_487, CLK, g465);
MUX2_X1 g_tmp_wire_488 (g4642, g465, SE, tmp_wire_488);
DFF_X1 g_g457 (tmp_wire_488, CLK, g457);
MUX2_X1 g_tmp_wire_489 (g6353, g457, SE, tmp_wire_489);
DFF_X1 g_g468 (tmp_wire_489, CLK, g468);
MUX2_X1 g_tmp_wire_490 (g4643, g468, SE, tmp_wire_490);
DFF_X1 g_g458 (tmp_wire_490, CLK, g458);
MUX2_X1 g_tmp_wire_491 (g6354, g458, SE, tmp_wire_491);
DFF_X1 g_g471 (tmp_wire_491, CLK, g471);
MUX2_X1 g_tmp_wire_492 (g4644, g471, SE, tmp_wire_492);
DFF_X1 g_g474 (tmp_wire_492, CLK, g474);
MUX2_X1 g_tmp_wire_493 (g6355, g474, SE, tmp_wire_493);
DFF_X1 g_g480 (tmp_wire_493, CLK, g480);
MUX2_X1 g_tmp_wire_494 (g4645, g480, SE, tmp_wire_494);
DFF_X1 g_g475 (tmp_wire_494, CLK, g475);
MUX2_X1 g_tmp_wire_495 (g6356, g475, SE, tmp_wire_495);
DFF_X1 g_g483 (tmp_wire_495, CLK, g483);
MUX2_X1 g_tmp_wire_496 (g4646, g483, SE, tmp_wire_496);
DFF_X1 g_g476 (tmp_wire_496, CLK, g476);
MUX2_X1 g_tmp_wire_497 (g6357, g476, SE, tmp_wire_497);
DFF_X1 g_g486 (tmp_wire_497, CLK, g486);
MUX2_X1 g_tmp_wire_498 (g4647, g486, SE, tmp_wire_498);
DFF_X1 g_g477 (tmp_wire_498, CLK, g477);
MUX2_X1 g_tmp_wire_499 (g6358, g477, SE, tmp_wire_499);
DFF_X1 g_g489 (tmp_wire_499, CLK, g489);
MUX2_X1 g_tmp_wire_500 (g4648, g489, SE, tmp_wire_500);
DFF_X1 g_g478 (tmp_wire_500, CLK, g478);
MUX2_X1 g_tmp_wire_501 (g6359, g478, SE, tmp_wire_501);
DFF_X1 g_g492 (tmp_wire_501, CLK, g492);
MUX2_X1 g_tmp_wire_502 (g4649, g492, SE, tmp_wire_502);
DFF_X1 g_g479 (tmp_wire_502, CLK, g479);
MUX2_X1 g_tmp_wire_503 (g6360, g479, SE, tmp_wire_503);
DFF_X1 g_g495 (tmp_wire_503, CLK, g495);
MUX2_X1 g_tmp_wire_504 (g4650, g495, SE, tmp_wire_504);
DFF_X1 g_g516 (tmp_wire_504, CLK, g516);
MUX2_X1 g_tmp_wire_505 (g6361, g516, SE, tmp_wire_505);
DFF_X1 g_g518 (tmp_wire_505, CLK, g518);
MUX2_X1 g_tmp_wire_506 (g4651, g518, SE, tmp_wire_506);
DFF_X1 g_g517 (tmp_wire_506, CLK, g517);
MUX2_X1 g_tmp_wire_507 (g6362, g517, SE, tmp_wire_507);
DFF_X1 g_g521 (tmp_wire_507, CLK, g521);
MUX2_X1 g_tmp_wire_508 (g3844, g521, SE, tmp_wire_508);
DFF_X1 g_g535 (tmp_wire_508, CLK, g535);
MUX2_X1 g_tmp_wire_509 (g6363, g535, SE, tmp_wire_509);
DFF_X1 g_g536 (tmp_wire_509, CLK, g536);
MUX2_X1 g_tmp_wire_510 (g3845, g536, SE, tmp_wire_510);
DFF_X1 g_g539 (tmp_wire_510, CLK, g539);
MUX2_X1 g_tmp_wire_511 (g6364, g539, SE, tmp_wire_511);
DFF_X1 g_g540 (tmp_wire_511, CLK, g540);
MUX2_X1 g_tmp_wire_512 (g3846, g540, SE, tmp_wire_512);
DFF_X1 g_g543 (tmp_wire_512, CLK, g543);
MUX2_X1 g_tmp_wire_513 (g6365, g543, SE, tmp_wire_513);
DFF_X1 g_g544 (tmp_wire_513, CLK, g544);
MUX2_X1 g_tmp_wire_514 (g9026, g544, SE, tmp_wire_514);
DFF_X1 g_g547 (tmp_wire_514, CLK, g547);
MUX2_X1 g_tmp_wire_515 (g9027, g547, SE, tmp_wire_515);
DFF_X1 g_g550 (tmp_wire_515, CLK, g550);
MUX2_X1 g_tmp_wire_516 (g9028, g550, SE, tmp_wire_516);
DFF_X1 g_g553 (tmp_wire_516, CLK, g553);
MUX2_X1 g_tmp_wire_517 (g3847, g553, SE, tmp_wire_517);
DFF_X1 g_g556 (tmp_wire_517, CLK, g556);
MUX2_X1 g_tmp_wire_518 (g6366, g556, SE, tmp_wire_518);
DFF_X1 g_g557 (tmp_wire_518, CLK, g557);
MUX2_X1 g_tmp_wire_519 (g3848, g557, SE, tmp_wire_519);
DFF_X1 g_g566 (tmp_wire_519, CLK, g566);
MUX2_X1 g_tmp_wire_520 (g6367, g566, SE, tmp_wire_520);
DFF_X1 g_g567 (tmp_wire_520, CLK, g567);
MUX2_X1 g_tmp_wire_521 (g3850, g567, SE, tmp_wire_521);
DFF_X1 g_g579 (tmp_wire_521, CLK, g579);
MUX2_X1 g_tmp_wire_522 (g6368, g579, SE, tmp_wire_522);
DFF_X1 g_g580 (tmp_wire_522, CLK, g580);
MUX2_X1 g_tmp_wire_523 (g3851, g580, SE, tmp_wire_523);
DFF_X1 g_g583 (tmp_wire_523, CLK, g583);
MUX2_X1 g_tmp_wire_524 (g6369, g583, SE, tmp_wire_524);
DFF_X1 g_g584 (tmp_wire_524, CLK, g584);
MUX2_X1 g_tmp_wire_525 (g3852, g584, SE, tmp_wire_525);
DFF_X1 g_g587 (tmp_wire_525, CLK, g587);
MUX2_X1 g_tmp_wire_526 (g6370, g587, SE, tmp_wire_526);
DFF_X1 g_g560 (tmp_wire_526, CLK, g560);
MUX2_X1 g_tmp_wire_527 (g9029, g560, SE, tmp_wire_527);
DFF_X1 g_g563 (tmp_wire_527, CLK, g563);
MUX2_X1 g_tmp_wire_528 (g9030, g563, SE, tmp_wire_528);
DFF_X1 g_g570 (tmp_wire_528, CLK, g570);
MUX2_X1 g_tmp_wire_529 (g9031, g570, SE, tmp_wire_529);
DFF_X1 g_g588 (tmp_wire_529, CLK, g588);
MUX2_X1 g_tmp_wire_530 (g9032, g588, SE, tmp_wire_530);
DFF_X1 g_g591 (tmp_wire_530, CLK, g591);
MUX2_X1 g_tmp_wire_531 (g9033, g591, SE, tmp_wire_531);
DFF_X1 g_g573 (tmp_wire_531, CLK, g573);
MUX2_X1 g_tmp_wire_532 (g3849, g573, SE, tmp_wire_532);
DFF_X1 g_g576 (tmp_wire_532, CLK, g576);
MUX2_X1 g_tmp_wire_533 (g576, g576, SE, tmp_wire_533);
DFF_X1 g_g595 (tmp_wire_533, CLK, g595);
MUX2_X1 g_tmp_wire_534 (g6795, g595, SE, tmp_wire_534);
DFF_X1 g_g596 (tmp_wire_534, CLK, g596);
MUX2_X1 g_tmp_wire_535 (g6796, g596, SE, tmp_wire_535);
DFF_X1 g_g597 (tmp_wire_535, CLK, g597);
MUX2_X1 g_tmp_wire_536 (g6797, g597, SE, tmp_wire_536);
DFF_X1 g_g598 (tmp_wire_536, CLK, g598);
MUX2_X1 g_tmp_wire_537 (g6798, g598, SE, tmp_wire_537);
DFF_X1 g_g599 (tmp_wire_537, CLK, g599);
MUX2_X1 g_tmp_wire_538 (g6807, g599, SE, tmp_wire_538);
DFF_X1 g_g600 (tmp_wire_538, CLK, g600);
MUX2_X1 g_tmp_wire_539 (g6799, g600, SE, tmp_wire_539);
DFF_X1 g_g601 (tmp_wire_539, CLK, g601);
MUX2_X1 g_tmp_wire_540 (g6800, g601, SE, tmp_wire_540);
DFF_X1 g_g602 (tmp_wire_540, CLK, g602);
MUX2_X1 g_tmp_wire_541 (g6801, g602, SE, tmp_wire_541);
DFF_X1 g_g603 (tmp_wire_541, CLK, g603);
MUX2_X1 g_tmp_wire_542 (g6802, g603, SE, tmp_wire_542);
DFF_X1 g_g604 (tmp_wire_542, CLK, g604);
MUX2_X1 g_tmp_wire_543 (g6803, g604, SE, tmp_wire_543);
DFF_X1 g_g605 (tmp_wire_543, CLK, g605);
MUX2_X1 g_tmp_wire_544 (g6804, g605, SE, tmp_wire_544);
DFF_X1 g_g606 (tmp_wire_544, CLK, g606);
MUX2_X1 g_tmp_wire_545 (g6805, g606, SE, tmp_wire_545);
DFF_X1 g_g607 (tmp_wire_545, CLK, g607);
MUX2_X1 g_tmp_wire_546 (g6806, g607, SE, tmp_wire_546);
DFF_X1 g_g608 (tmp_wire_546, CLK, g608);
MUX2_X1 g_tmp_wire_547 (g6808, g608, SE, tmp_wire_547);
DFF_X1 g_g609 (tmp_wire_547, CLK, g609);
MUX2_X1 g_tmp_wire_548 (g6809, g609, SE, tmp_wire_548);
DFF_X1 g_g610 (tmp_wire_548, CLK, g610);
MUX2_X1 g_tmp_wire_549 (g6810, g610, SE, tmp_wire_549);
DFF_X1 g_g611 (tmp_wire_549, CLK, g611);
MUX2_X1 g_tmp_wire_550 (g6811, g611, SE, tmp_wire_550);
DFF_X1 g_g612 (tmp_wire_550, CLK, g612);
MUX2_X1 g_tmp_wire_551 (g6820, g612, SE, tmp_wire_551);
DFF_X1 g_g613 (tmp_wire_551, CLK, g613);
MUX2_X1 g_tmp_wire_552 (g6812, g613, SE, tmp_wire_552);
DFF_X1 g_g614 (tmp_wire_552, CLK, g614);
MUX2_X1 g_tmp_wire_553 (g6813, g614, SE, tmp_wire_553);
DFF_X1 g_g615 (tmp_wire_553, CLK, g615);
MUX2_X1 g_tmp_wire_554 (g6814, g615, SE, tmp_wire_554);
DFF_X1 g_g616 (tmp_wire_554, CLK, g616);
MUX2_X1 g_tmp_wire_555 (g6815, g616, SE, tmp_wire_555);
DFF_X1 g_g617 (tmp_wire_555, CLK, g617);
MUX2_X1 g_tmp_wire_556 (g6816, g617, SE, tmp_wire_556);
DFF_X1 g_g618 (tmp_wire_556, CLK, g618);
MUX2_X1 g_tmp_wire_557 (g6817, g618, SE, tmp_wire_557);
DFF_X1 g_g619 (tmp_wire_557, CLK, g619);
MUX2_X1 g_tmp_wire_558 (g6818, g619, SE, tmp_wire_558);
DFF_X1 g_g620 (tmp_wire_558, CLK, g620);
MUX2_X1 g_tmp_wire_559 (g6819, g620, SE, tmp_wire_559);
DFF_X1 g_g621 (tmp_wire_559, CLK, g621);
MUX2_X1 g_tmp_wire_560 (g6821, g621, SE, tmp_wire_560);
DFF_X1 g_g622 (tmp_wire_560, CLK, g622);
MUX2_X1 g_tmp_wire_561 (g6822, g622, SE, tmp_wire_561);
DFF_X1 g_g623 (tmp_wire_561, CLK, g623);
MUX2_X1 g_tmp_wire_562 (g6831, g623, SE, tmp_wire_562);
DFF_X1 g_g624 (tmp_wire_562, CLK, g624);
MUX2_X1 g_tmp_wire_563 (g6823, g624, SE, tmp_wire_563);
DFF_X1 g_g625 (tmp_wire_563, CLK, g625);
MUX2_X1 g_tmp_wire_564 (g6824, g625, SE, tmp_wire_564);
DFF_X1 g_g626 (tmp_wire_564, CLK, g626);
MUX2_X1 g_tmp_wire_565 (g6825, g626, SE, tmp_wire_565);
DFF_X1 g_g627 (tmp_wire_565, CLK, g627);
MUX2_X1 g_tmp_wire_566 (g6826, g627, SE, tmp_wire_566);
DFF_X1 g_g628 (tmp_wire_566, CLK, g628);
MUX2_X1 g_tmp_wire_567 (g6827, g628, SE, tmp_wire_567);
DFF_X1 g_g629 (tmp_wire_567, CLK, g629);
MUX2_X1 g_tmp_wire_568 (g6828, g629, SE, tmp_wire_568);
DFF_X1 g_g630 (tmp_wire_568, CLK, g630);
MUX2_X1 g_tmp_wire_569 (g6829, g630, SE, tmp_wire_569);
DFF_X1 g_g631 (tmp_wire_569, CLK, g631);
MUX2_X1 g_tmp_wire_570 (g6830, g631, SE, tmp_wire_570);
DFF_X1 g_g632 (tmp_wire_570, CLK, g632);
MUX2_X1 g_tmp_wire_571 (g4652, g632, SE, tmp_wire_571);
DFF_X1 g_g646 (tmp_wire_571, CLK, g646);
MUX2_X1 g_tmp_wire_572 (g646, g646, SE, tmp_wire_572);
DFF_X1 g_g652 (tmp_wire_572, CLK, g652);
MUX2_X1 g_tmp_wire_573 (g7743, g652, SE, tmp_wire_573);
DFF_X1 g_g661 (tmp_wire_573, CLK, g661);
MUX2_X1 g_tmp_wire_574 (g7744, g661, SE, tmp_wire_574);
DFF_X1 g_g665 (tmp_wire_574, CLK, g665);
MUX2_X1 g_tmp_wire_575 (g7745, g665, SE, tmp_wire_575);
DFF_X1 g_g669 (tmp_wire_575, CLK, g669);
MUX2_X1 g_tmp_wire_576 (g7746, g669, SE, tmp_wire_576);
DFF_X1 g_g673 (tmp_wire_576, CLK, g673);
MUX2_X1 g_tmp_wire_577 (g7747, g673, SE, tmp_wire_577);
DFF_X1 g_g677 (tmp_wire_577, CLK, g677);
MUX2_X1 g_tmp_wire_578 (g7748, g677, SE, tmp_wire_578);
DFF_X1 g_g681 (tmp_wire_578, CLK, g681);
MUX2_X1 g_tmp_wire_579 (g7749, g681, SE, tmp_wire_579);
DFF_X1 g_g685 (tmp_wire_579, CLK, g685);
MUX2_X1 g_tmp_wire_580 (g7750, g685, SE, tmp_wire_580);
DFF_X1 g_g706 (tmp_wire_580, CLK, g706);
MUX2_X1 g_tmp_wire_581 (g7751, g706, SE, tmp_wire_581);
DFF_X1 g_g710 (tmp_wire_581, CLK, g710);
MUX2_X1 g_tmp_wire_582 (g7752, g710, SE, tmp_wire_582);
DFF_X1 g_g714 (tmp_wire_582, CLK, g714);
MUX2_X1 g_tmp_wire_583 (g7753, g714, SE, tmp_wire_583);
DFF_X1 g_g718 (tmp_wire_583, CLK, g718);
MUX2_X1 g_tmp_wire_584 (g7755, g718, SE, tmp_wire_584);
DFF_X1 g_g734 (tmp_wire_584, CLK, g734);
MUX2_X1 g_tmp_wire_585 (g7754, g734, SE, tmp_wire_585);
DFF_X1 g_g730 (tmp_wire_585, CLK, g730);
MUX2_X1 g_tmp_wire_586 (g6371, g730, SE, tmp_wire_586);
DFF_X1 g_g689 (tmp_wire_586, CLK, g689);
MUX2_X1 g_tmp_wire_587 (g6840, g689, SE, tmp_wire_587);
DFF_X1 g_g758 (tmp_wire_587, CLK, g758);
MUX2_X1 g_tmp_wire_588 (g6832, g758, SE, tmp_wire_588);
DFF_X1 g_g759 (tmp_wire_588, CLK, g759);
MUX2_X1 g_tmp_wire_589 (g6833, g759, SE, tmp_wire_589);
DFF_X1 g_g760 (tmp_wire_589, CLK, g760);
MUX2_X1 g_tmp_wire_590 (g6834, g760, SE, tmp_wire_590);
DFF_X1 g_g761 (tmp_wire_590, CLK, g761);
MUX2_X1 g_tmp_wire_591 (g6835, g761, SE, tmp_wire_591);
DFF_X1 g_g762 (tmp_wire_591, CLK, g762);
MUX2_X1 g_tmp_wire_592 (g6836, g762, SE, tmp_wire_592);
DFF_X1 g_g763 (tmp_wire_592, CLK, g763);
MUX2_X1 g_tmp_wire_593 (g6837, g763, SE, tmp_wire_593);
DFF_X1 g_g764 (tmp_wire_593, CLK, g764);
MUX2_X1 g_tmp_wire_594 (g6838, g764, SE, tmp_wire_594);
DFF_X1 g_g765 (tmp_wire_594, CLK, g765);
MUX2_X1 g_tmp_wire_595 (g6839, g765, SE, tmp_wire_595);
DFF_X1 g_g766 (tmp_wire_595, CLK, g766);
MUX2_X1 g_tmp_wire_596 (g6841, g766, SE, tmp_wire_596);
DFF_X1 g_g767 (tmp_wire_596, CLK, g767);
MUX2_X1 g_tmp_wire_597 (g6842, g767, SE, tmp_wire_597);
DFF_X1 g_g768 (tmp_wire_597, CLK, g768);
MUX2_X1 g_tmp_wire_598 (g6843, g768, SE, tmp_wire_598);
DFF_X1 g_g769 (tmp_wire_598, CLK, g769);
MUX2_X1 g_tmp_wire_599 (g6844, g769, SE, tmp_wire_599);
DFF_X1 g_g770 (tmp_wire_599, CLK, g770);
MUX2_X1 g_tmp_wire_600 (g6845, g770, SE, tmp_wire_600);
DFF_X1 g_g771 (tmp_wire_600, CLK, g771);
MUX2_X1 g_tmp_wire_601 (g6846, g771, SE, tmp_wire_601);
DFF_X1 g_g772 (tmp_wire_601, CLK, g772);
MUX2_X1 g_tmp_wire_602 (g6847, g772, SE, tmp_wire_602);
DFF_X1 g_g773 (tmp_wire_602, CLK, g773);
MUX2_X1 g_tmp_wire_603 (g6848, g773, SE, tmp_wire_603);
DFF_X1 g_g774 (tmp_wire_603, CLK, g774);
MUX2_X1 g_tmp_wire_604 (g3854, g774, SE, tmp_wire_604);
DFF_X1 g_g795 (tmp_wire_604, CLK, g795);
MUX2_X1 g_tmp_wire_605 (g5162, g795, SE, tmp_wire_605);
DFF_X1 g_g792 (tmp_wire_605, CLK, g792);
MUX2_X1 g_tmp_wire_606 (g5734, g792, SE, tmp_wire_606);
DFF_X1 g_g782 (tmp_wire_606, CLK, g782);
MUX2_X1 g_tmp_wire_607 (g7756, g782, SE, tmp_wire_607);
DFF_X1 g_g799 (tmp_wire_607, CLK, g799);
MUX2_X1 g_tmp_wire_608 (g7757, g799, SE, tmp_wire_608);
DFF_X1 g_g803 (tmp_wire_608, CLK, g803);
MUX2_X1 g_tmp_wire_609 (g7510, g803, SE, tmp_wire_609);
DFF_X1 g_g806 (tmp_wire_609, CLK, g806);
MUX2_X1 g_tmp_wire_610 (g7511, g806, SE, tmp_wire_610);
DFF_X1 g_g809 (tmp_wire_610, CLK, g809);
MUX2_X1 g_tmp_wire_611 (g7758, g809, SE, tmp_wire_611);
DFF_X1 g_g812 (tmp_wire_611, CLK, g812);
MUX2_X1 g_tmp_wire_612 (g7759, g812, SE, tmp_wire_612);
DFF_X1 g_g775 (tmp_wire_612, CLK, g775);
MUX2_X1 g_tmp_wire_613 (g7296, g775, SE, tmp_wire_613);
DFF_X1 g_g778 (tmp_wire_613, CLK, g778);
MUX2_X1 g_tmp_wire_614 (g7760, g778, SE, tmp_wire_614);
DFF_X1 g_g815 (tmp_wire_614, CLK, g815);
MUX2_X1 g_tmp_wire_615 (g7761, g815, SE, tmp_wire_615);
DFF_X1 g_g819 (tmp_wire_615, CLK, g819);
MUX2_X1 g_tmp_wire_616 (g7512, g819, SE, tmp_wire_616);
DFF_X1 g_g822 (tmp_wire_616, CLK, g822);
MUX2_X1 g_tmp_wire_617 (g7513, g822, SE, tmp_wire_617);
DFF_X1 g_g825 (tmp_wire_617, CLK, g825);
MUX2_X1 g_tmp_wire_618 (g7762, g825, SE, tmp_wire_618);
DFF_X1 g_g828 (tmp_wire_618, CLK, g828);
MUX2_X1 g_tmp_wire_619 (g7763, g828, SE, tmp_wire_619);
DFF_X1 g_g786 (tmp_wire_619, CLK, g786);
MUX2_X1 g_tmp_wire_620 (g7297, g786, SE, tmp_wire_620);
DFF_X1 g_g789 (tmp_wire_620, CLK, g789);
MUX2_X1 g_tmp_wire_621 (g3857, g789, SE, tmp_wire_621);
DFF_X1 g_g955 (tmp_wire_621, CLK, g955);
MUX2_X1 g_tmp_wire_622 (g5169, g955, SE, tmp_wire_622);
DFF_X1 g_g959 (tmp_wire_622, CLK, g959);
MUX2_X1 g_tmp_wire_623 (g5170, g959, SE, tmp_wire_623);
DFF_X1 g_g945 (tmp_wire_623, CLK, g945);
MUX2_X1 g_tmp_wire_624 (g8664, g945, SE, tmp_wire_624);
DFF_X1 g_g948 (tmp_wire_624, CLK, g948);
MUX2_X1 g_tmp_wire_625 (g8665, g948, SE, tmp_wire_625);
DFF_X1 g_g949 (tmp_wire_625, CLK, g949);
MUX2_X1 g_tmp_wire_626 (g8666, g949, SE, tmp_wire_626);
DFF_X1 g_g950 (tmp_wire_626, CLK, g950);
MUX2_X1 g_tmp_wire_627 (g8667, g950, SE, tmp_wire_627);
DFF_X1 g_g951 (tmp_wire_627, CLK, g951);
MUX2_X1 g_tmp_wire_628 (g8668, g951, SE, tmp_wire_628);
DFF_X1 g_g952 (tmp_wire_628, CLK, g952);
MUX2_X1 g_tmp_wire_629 (g8669, g952, SE, tmp_wire_629);
DFF_X1 g_g953 (tmp_wire_629, CLK, g953);
MUX2_X1 g_tmp_wire_630 (g8670, g953, SE, tmp_wire_630);
DFF_X1 g_g954 (tmp_wire_630, CLK, g954);
MUX2_X1 g_tmp_wire_631 (g8671, g954, SE, tmp_wire_631);
DFF_X1 g_g943 (tmp_wire_631, CLK, g943);
MUX2_X1 g_tmp_wire_632 (g5168, g943, SE, tmp_wire_632);
DFF_X1 g_g936 (tmp_wire_632, CLK, g936);
MUX2_X1 g_tmp_wire_633 (g5735, g936, SE, tmp_wire_633);
DFF_X1 g_g940 (tmp_wire_633, CLK, g940);
MUX2_X1 g_tmp_wire_634 (g2652, g940, SE, tmp_wire_634);
DFF_X1 g_g942 (tmp_wire_634, CLK, g942);
MUX2_X1 g_tmp_wire_635 (g6372, g942, SE, tmp_wire_635);
DFF_X1 g_g944 (tmp_wire_635, CLK, g944);
MUX2_X1 g_tmp_wire_636 (g8220, g944, SE, tmp_wire_636);
DFF_X1 g_g855 (tmp_wire_636, CLK, g855);
MUX2_X1 g_tmp_wire_637 (g8221, g855, SE, tmp_wire_637);
DFF_X1 g_g859 (tmp_wire_637, CLK, g859);
MUX2_X1 g_tmp_wire_638 (g8222, g859, SE, tmp_wire_638);
DFF_X1 g_g863 (tmp_wire_638, CLK, g863);
MUX2_X1 g_tmp_wire_639 (g2651, g863, SE, tmp_wire_639);
DFF_X1 g_g831 (tmp_wire_639, CLK, g831);
MUX2_X1 g_tmp_wire_640 (g2650, g831, SE, tmp_wire_640);
DFF_X1 g_g834 (tmp_wire_640, CLK, g834);
MUX2_X1 g_tmp_wire_641 (g2649, g834, SE, tmp_wire_641);
DFF_X1 g_g837 (tmp_wire_641, CLK, g837);
MUX2_X1 g_tmp_wire_642 (g2648, g837, SE, tmp_wire_642);
DFF_X1 g_g840 (tmp_wire_642, CLK, g840);
MUX2_X1 g_tmp_wire_643 (g2647, g840, SE, tmp_wire_643);
DFF_X1 g_g843 (tmp_wire_643, CLK, g843);
MUX2_X1 g_tmp_wire_644 (g2646, g843, SE, tmp_wire_644);
DFF_X1 g_g846 (tmp_wire_644, CLK, g846);
MUX2_X1 g_tmp_wire_645 (g2645, g846, SE, tmp_wire_645);
DFF_X1 g_g849 (tmp_wire_645, CLK, g849);
MUX2_X1 g_tmp_wire_646 (g2644, g849, SE, tmp_wire_646);
DFF_X1 g_g852 (tmp_wire_646, CLK, g852);
MUX2_X1 g_tmp_wire_647 (g7102, g852, SE, tmp_wire_647);
DFF_X1 g_g890 (tmp_wire_647, CLK, g890);
MUX2_X1 g_tmp_wire_648 (g890, g890, SE, tmp_wire_648);
DFF_X1 g_g878 (tmp_wire_648, CLK, g878);
MUX2_X1 g_tmp_wire_649 (g878, g878, SE, tmp_wire_649);
DFF_X1 g_g926 (tmp_wire_649, CLK, g926);
MUX2_X1 g_tmp_wire_650 (g5165, g926, SE, tmp_wire_650);
DFF_X1 g_g875 (tmp_wire_650, CLK, g875);
MUX2_X1 g_tmp_wire_651 (g5163, g875, SE, tmp_wire_651);
DFF_X1 g_g866 (tmp_wire_651, CLK, g866);
MUX2_X1 g_tmp_wire_652 (g3856, g866, SE, tmp_wire_652);
DFF_X1 g_g929 (tmp_wire_652, CLK, g929);
MUX2_X1 g_tmp_wire_653 (g5166, g929, SE, tmp_wire_653);
DFF_X1 g_g933 (tmp_wire_653, CLK, g933);
MUX2_X1 g_tmp_wire_654 (g5167, g933, SE, tmp_wire_654);
DFF_X1 g_g871 (tmp_wire_654, CLK, g871);
MUX2_X1 g_tmp_wire_655 (g4654, g871, SE, tmp_wire_655);
DFF_X1 g_g874 (tmp_wire_655, CLK, g874);
MUX2_X1 g_tmp_wire_656 (g3855, g874, SE, tmp_wire_656);
DFF_X1 g_g891 (tmp_wire_656, CLK, g891);
MUX2_X1 g_tmp_wire_657 (g891, g891, SE, tmp_wire_657);
DFF_X1 g_g896 (tmp_wire_657, CLK, g896);
MUX2_X1 g_tmp_wire_658 (g896, g896, SE, tmp_wire_658);
DFF_X1 g_g901 (tmp_wire_658, CLK, g901);
MUX2_X1 g_tmp_wire_659 (g901, g901, SE, tmp_wire_659);
DFF_X1 g_g906 (tmp_wire_659, CLK, g906);
MUX2_X1 g_tmp_wire_660 (g906, g906, SE, tmp_wire_660);
DFF_X1 g_g911 (tmp_wire_660, CLK, g911);
MUX2_X1 g_tmp_wire_661 (g911, g911, SE, tmp_wire_661);
DFF_X1 g_g916 (tmp_wire_661, CLK, g916);
MUX2_X1 g_tmp_wire_662 (g916, g916, SE, tmp_wire_662);
DFF_X1 g_g921 (tmp_wire_662, CLK, g921);
MUX2_X1 g_tmp_wire_663 (g921, g921, SE, tmp_wire_663);
DFF_X1 g_g883 (tmp_wire_663, CLK, g883);
MUX2_X1 g_tmp_wire_664 (g7099, g883, SE, tmp_wire_664);
DFF_X1 g_g887 (tmp_wire_664, CLK, g887);
MUX2_X1 g_tmp_wire_665 (g7100, g887, SE, tmp_wire_665);
DFF_X1 g_g888 (tmp_wire_665, CLK, g888);
MUX2_X1 g_tmp_wire_666 (g7101, g888, SE, tmp_wire_666);
DFF_X1 g_g889 (tmp_wire_666, CLK, g889);
MUX2_X1 g_tmp_wire_667 (g9386, g889, SE, tmp_wire_667);
DFF_X1 g_g741 (tmp_wire_667, CLK, g741);
MUX2_X1 g_tmp_wire_668 (g8956, g741, SE, tmp_wire_668);
DFF_X1 g_g746 (tmp_wire_668, CLK, g746);
BUF_X1 g_SO (g746, SO);
INV_X1 g_I5353 (g3833, I5353);
INV_X1 g_g206 (I5353, g206);
INV_X1 g_I5356 (g3837, I5356);
INV_X1 g_g291 (I5356, g291);
INV_X1 g_I5359 (g3839, I5359);
INV_X1 g_g372 (I5359, g372);
INV_X1 g_I5362 (g3841, I5362);
INV_X1 g_g453 (I5362, g453);
INV_X1 g_I5365 (g3843, I5365);
INV_X1 g_g534 (I5365, g534);
INV_X1 g_I5368 (g3853, I5368);
INV_X1 g_g594 (I5368, g594);
INV_X1 g_I5371 (g633, I5371);
INV_X1 g_g636 (I5371, g636);
INV_X1 g_I5374 (g634, I5374);
INV_X1 g_g639 (I5374, g639);
INV_X1 g_I5377 (g635, I5377);
INV_X1 g_g642 (I5377, g642);
INV_X1 g_I5380 (g645, I5380);
INV_X1 g_g649 (I5380, g649);
INV_X1 g_I5383 (g647, I5383);
INV_X1 g_g655 (I5383, g655);
INV_X1 g_I5386 (g648, I5386);
INV_X1 g_g658 (I5386, g658);
INV_X1 g_I5389 (g690, I5389);
INV_X1 g_g691 (I5389, g691);
INV_X1 g_I5392 (g694, I5392);
INV_X1 g_g695 (I5392, g695);
INV_X1 g_I5395 (g698, I5395);
INV_X1 g_g699 (I5395, g699);
INV_X1 g_I5398 (g702, I5398);
INV_X1 g_g703 (I5398, g703);
INV_X1 g_I5401 (g723, I5401);
INV_X1 g_g724 (I5401, g724);
INV_X1 g_I5404 (g722, I5404);
INV_X1 g_g738 (I5404, g738);
INV_X1 g_I5407 (g4653, I5407);
INV_X1 g_g785 (I5407, g785);
INV_X1 g_I5410 (g8866, I5410);
INV_X1 g_g1006 (I5410, g1006);
INV_X1 g_I5413 (g1016, I5413);
INV_X1 g_g1011 (I5413, g1011);
INV_X1 g_I5416 (g8868, I5416);
INV_X1 g_g1015 (I5416, g1015);
INV_X1 g_I5419 (g1603, I5419);
INV_X1 g_g1017 (I5419, g1017);
INV_X1 g_I5422 (g1234, I5422);
INV_X1 g_g1235 (I5422, g1235);
INV_X1 g_I5425 (g1245, I5425);
INV_X1 g_g1246 (I5425, g1246);
INV_X1 g_I5428 (g49, I5428);
INV_X1 g_g1555 (I5428, g1555);
INV_X1 g_g1556 (g65, g1556);
INV_X1 g_I5432 (g1176, I5432);
INV_X1 g_g1557 (I5432, g1557);
INV_X1 g_I5435 (g1461, I5435);
INV_X1 g_g1558 (I5435, g1558);
INV_X1 g_g1562 (g636, g1562);
INV_X1 g_g1563 (g639, g1563);
INV_X1 g_g1564 (g642, g1564);
INV_X1 g_g1565 (g649, g1565);
INV_X1 g_g1566 (g652, g1566);
INV_X1 g_g1567 (g655, g1567);
INV_X1 g_g1568 (g658, g1568);
INV_X1 g_g1569 (g661, g1569);
INV_X1 g_g1570 (g665, g1570);
INV_X1 g_g1571 (g669, g1571);
INV_X1 g_g1572 (g673, g1572);
INV_X1 g_g1573 (g677, g1573);
INV_X1 g_g1574 (g681, g1574);
INV_X1 g_g1575 (g685, g1575);
INV_X1 g_g1576 (g691, g1576);
INV_X1 g_g1577 (g695, g1577);
INV_X1 g_g1578 (g699, g1578);
INV_X1 g_g1579 (g703, g1579);
INV_X1 g_g1580 (g706, g1580);
INV_X1 g_g1581 (g710, g1581);
INV_X1 g_g1582 (g714, g1582);
INV_X1 g_g1583 (g718, g1583);
INV_X1 g_g1584 (g738, g1584);
INV_X1 g_g1585 (g724, g1585);
INV_X1 g_g1586 (g730, g1586);
INV_X1 g_g1587 (g734, g1587);
INV_X1 g_g1588 (g741, g1588);
INV_X1 g_g1589 (g746, g1589);
INV_X1 g_I5466 (g926, I5466);
INV_X1 g_g1590 (I5466, g1590);
INV_X1 g_g1597 (g973, g1597);
INV_X1 g_g1600 (g976, g1600);
INV_X1 g_I5471 (g1029, I5471);
INV_X1 g_g1603 (I5471, g1603);
INV_X1 g_g1611 (g1073, g1611);
INV_X1 g_I5475 (g1084, I5475);
INV_X1 g_g1612 (I5475, g1612);
INV_X1 g_I5478 (g1148, I5478);
INV_X1 g_g1616 (I5478, g1616);
INV_X1 g_g1637 (g1087, g1637);
INV_X1 g_g1638 (g1092, g1638);
INV_X1 g_g1639 (g1207, g1639);
INV_X1 g_g1643 (g1211, g1643);
INV_X1 g_g1646 (g1214, g1646);
INV_X1 g_g1649 (g1217, g1649);
INV_X1 g_g1652 (g1220, g1652);
INV_X1 g_g1655 (g1231, g1655);
INV_X1 g_g1658 (g1313, g1658);
INV_X1 g_g1661 (g1405, g1661);
INV_X1 g_g1662 (g1412, g1662);
INV_X1 g_g1663 (g1416, g1663);
INV_X1 g_g1664 (g1462, g1664);
INV_X1 g_g1665 (g1467, g1665);
INV_X1 g_g1666 (g1472, g1666);
INV_X1 g_g1667 (g1481, g1667);
INV_X1 g_g1670 (g1489, g1670);
INV_X1 g_g1671 (g1494, g1671);
INV_X1 g_g1672 (g1499, g1672);
INV_X1 g_g1673 (g1504, g1673);
INV_X1 g_g1674 (g1514, g1674);
INV_X1 g_g1675 (g1519, g1675);
INV_X1 g_g1676 (g727, g1676);
INV_X1 g_g1677 (g1532, g1677);
INV_X1 g_I5512 (g557, I5512);
INV_X1 g_g1679 (I5512, g1679);
INV_X1 g_I5515 (g567, I5515);
INV_X1 g_g1680 (I5515, g1680);
INV_X1 g_g1681 (g929, g1681);
INV_X1 g_g1683 (g795, g1683);
INV_X1 g_g1684 (g1, g1684);
INV_X1 g_I5528 (g43, I5528);
INV_X1 g_g1685 (I5528, g1685);
INV_X1 g_I5531 (g866, I5531);
INV_X1 g_g1686 (I5531, g1686);
INV_X1 g_g1687 (g10, g1687);
INV_X1 g_I5535 (g48, I5535);
INV_X1 g_g1688 (I5535, g1688);
INV_X1 g_g1689 (g855, g1689);
INV_X1 g_g1694 (g21, g1694);
INV_X1 g_g1695 (g778, g1695);
INV_X1 g_I5542 (g1272, I5542);
INV_X1 g_g1698 (I5542, g1698);
INV_X1 g_I5545 (g1276, I5545);
INV_X1 g_g1701 (I5545, g1701);
INV_X1 g_I5548 (g1280, I5548);
INV_X1 g_g1704 (I5548, g1704);
INV_X1 g_g1707 (g955, g1707);
INV_X1 g_I5552 (g1284, I5552);
INV_X1 g_g1708 (I5552, g1708);
INV_X1 g_I5555 (g1288, I5555);
INV_X1 g_g1711 (I5555, g1711);
INV_X1 g_I5559 (g1292, I5559);
INV_X1 g_g1715 (I5559, g1715);
INV_X1 g_I5562 (g1300, I5562);
INV_X1 g_g1718 (I5562, g1718);
INV_X1 g_I5565 (g1296, I5565);
INV_X1 g_g1721 (I5565, g1721);
INV_X1 g_I5568 (g1409, I5568);
INV_X1 g_g1724 (I5568, g1724);
INV_X1 g_g1726 (g158, g1726);
INV_X1 g_g1727 (g596, g1727);
INV_X1 g_g1732 (g1439, g1732);
INV_X1 g_I5577 (g172, I5577);
INV_X1 g_g1736 (I5577, g1736);
INV_X1 g_g1737 (g597, g1737);
INV_X1 g_g1738 (g741, g1738);
INV_X1 g_g1742 (g1486, g1742);
INV_X1 g_g1743 (g598, g1743);
INV_X1 g_g1744 (g600, g1744);
INV_X1 g_g1745 (g746, g1745);
INV_X1 g_g1746 (g290, g1746);
INV_X1 g_g1747 (g599, g1747);
INV_X1 g_g1748 (g601, g1748);
INV_X1 g_g1749 (g371, g1749);
INV_X1 g_g1750 (g602, g1750);
INV_X1 g_g1751 (g452, g1751);
INV_X1 g_g1752 (g603, g1752);
INV_X1 g_g1756 (g533, g1756);
INV_X1 g_g1757 (g604, g1757);
INV_X1 g_g1758 (g1084, g1758);
INV_X1 g_I5605 (g58, I5605);
INV_X1 g_g1760 (I5605, g1760);
INV_X1 g_g1768 (g605, g1768);
INV_X1 g_I5609 (g16, I5609);
INV_X1 g_g1769 (I5609, g1769);
INV_X1 g_g1770 (g606, g1770);
INV_X1 g_g1771 (g609, g1771);
INV_X1 g_g1772 (g607, g1772);
INV_X1 g_g1773 (g610, g1773);
INV_X1 g_I5616 (g979, I5616);
INV_X1 g_g1774 (I5616, g1774);
INV_X1 g_g1776 (g608, g1776);
INV_X1 g_g1777 (g611, g1777);
INV_X1 g_g1778 (g613, g1778);
INV_X1 g_g1779 (g612, g1779);
INV_X1 g_g1780 (g614, g1780);
INV_X1 g_g1781 (g622, g1781);
INV_X1 g_g1782 (g624, g1782);
INV_X1 g_I5633 (g891, I5633);
INV_X1 g_g1783 (I5633, g1783);
INV_X1 g_I5636 (g891, I5636);
INV_X1 g_g1784 (I5636, g1784);
INV_X1 g_g1785 (g615, g1785);
INV_X1 g_g1786 (g623, g1786);
INV_X1 g_g1787 (g625, g1787);
INV_X1 g_g1788 (g984, g1788);
INV_X1 g_g1789 (g1034, g1789);
INV_X1 g_g1792 (g616, g1792);
INV_X1 g_g1793 (g626, g1793);
INV_X1 g_I5646 (g883, I5646);
INV_X1 g_g1794 (I5646, g1794);
INV_X1 g_I5649 (g1389, I5649);
INV_X1 g_g1795 (I5649, g1795);
INV_X1 g_g1796 (g617, g1796);
INV_X1 g_g1797 (g627, g1797);
INV_X1 g_I5654 (g921, I5654);
INV_X1 g_g1798 (I5654, g1798);
INV_X1 g_I5657 (g921, I5657);
INV_X1 g_g1799 (I5657, g1799);
INV_X1 g_g1800 (g1477, g1800);
INV_X1 g_g1801 (g618, g1801);
INV_X1 g_g1802 (g628, g1802);
INV_X1 g_g1803 (g758, g1803);
INV_X1 g_I5664 (g916, I5664);
INV_X1 g_g1804 (I5664, g1804);
INV_X1 g_I5667 (g916, I5667);
INV_X1 g_g1805 (I5667, g1805);
INV_X1 g_I5670 (g941, I5670);
INV_X1 g_g1806 (I5670, g1806);
INV_X1 g_g1807 (g619, g1807);
INV_X1 g_g1808 (g629, g1808);
INV_X1 g_g1809 (g759, g1809);
INV_X1 g_I5676 (g911, I5676);
INV_X1 g_g1810 (I5676, g1810);
INV_X1 g_I5679 (g911, I5679);
INV_X1 g_g1811 (I5679, g1811);
INV_X1 g_I5682 (g168, I5682);
INV_X1 g_g1812 (I5682, g1812);
INV_X1 g_g1813 (g620, g1813);
INV_X1 g_g1814 (g630, g1814);
INV_X1 g_g1815 (g760, g1815);
INV_X1 g_g1816 (g767, g1816);
INV_X1 g_I5689 (g906, I5689);
INV_X1 g_g1817 (I5689, g1817);
INV_X1 g_I5692 (g906, I5692);
INV_X1 g_g1818 (I5692, g1818);
INV_X1 g_g1820 (g621, g1820);
INV_X1 g_g1821 (g631, g1821);
INV_X1 g_g1822 (g761, g1822);
INV_X1 g_g1823 (g768, g1823);
INV_X1 g_I5706 (g901, I5706);
INV_X1 g_g1824 (I5706, g1824);
INV_X1 g_I5709 (g901, I5709);
INV_X1 g_g1825 (I5709, g1825);
INV_X1 g_g1826 (g632, g1826);
INV_X1 g_g1827 (g762, g1827);
INV_X1 g_g1828 (g769, g1828);
INV_X1 g_I5715 (g896, I5715);
INV_X1 g_g1829 (I5715, g1829);
INV_X1 g_I5718 (g896, I5718);
INV_X1 g_g1830 (I5718, g1830);
INV_X1 g_g1831 (g689, g1831);
INV_X1 g_g1832 (g763, g1832);
INV_X1 g_g1833 (g770, g1833);
INV_X1 g_g1837 (g1007, g1837);
INV_X1 g_g1838 (g1450, g1838);
INV_X1 g_g1842 (g764, g1842);
INV_X1 g_g1843 (g771, g1843);
INV_X1 g_g1847 (g765, g1847);
INV_X1 g_g1848 (g772, g1848);
INV_X1 g_I5732 (g859, I5732);
INV_X1 g_g1849 (I5732, g1849);
INV_X1 g_g1852 (g887, g1852);
INV_X1 g_g1853 (g766, g1853);
INV_X1 g_g1854 (g773, g1854);
INV_X1 g_g1855 (g866, g1855);
INV_X1 g_g1856 (g774, g1856);
INV_X1 g_g1857 (g889, g1857);
INV_X1 g_g1860 (g162, g1860);
INV_X1 g_g1863 (g68, g1863);
INV_X1 g_g1864 (g162, g1864);
INV_X1 g_g1865 (g1013, g1865);
INV_X1 g_g1866 (g71, g1866);
INV_X1 g_g1867 (g878, g1867);
INV_X1 g_I5747 (g1260, I5747);
INV_X1 g_g1868 (I5747, g1868);
INV_X1 g_g1869 (g74, g1869);
INV_X1 g_I5751 (g963, I5751);
INV_X1 g_g1870 (I5751, g1870);
INV_X1 g_I5754 (g966, I5754);
INV_X1 g_g1871 (I5754, g1871);
INV_X1 g_g1876 (g77, g1876);
INV_X1 g_g1877 (g595, g1877);
INV_X1 g_g1878 (g80, g1878);
INV_X1 g_I5763 (g1207, I5763);
INV_X1 g_g1879 (I5763, g1879);
INV_X1 g_I5766 (g1254, I5766);
INV_X1 g_g1886 (I5766, g1886);
INV_X1 g_g1887 (g83, g1887);
INV_X1 g_g1888 (g781, g1888);
INV_X1 g_g1889 (g1018, g1889);
INV_X1 g_I5772 (g1240, I5772);
INV_X1 g_g1894 (I5772, g1894);
INV_X1 g_I5775 (g1240, I5775);
INV_X1 g_g1895 (I5775, g1895);
INV_X1 g_g1896 (g86, g1896);
INV_X1 g_g1897 (g789, g1897);
INV_X1 g_I5781 (g979, I5781);
INV_X1 g_g1901 (I5781, g1901);
INV_X1 g_g1904 (g1021, g1904);
INV_X1 g_g1907 (g52, g1907);
INV_X1 g_g1908 (g812, g1908);
INV_X1 g_g1909 (g998, g1909);
INV_X1 g_I5789 (g1524, I5789);
INV_X1 g_g1911 (I5789, g1911);
INV_X1 g_g1912 (g1524, g1912);
INV_X1 g_g1916 (g775, g1916);
INV_X1 g_I5795 (g1236, I5795);
INV_X1 g_g1917 (I5795, g1917);
INV_X1 g_g1918 (g822, g1918);
INV_X1 g_g1922 (g1251, g1922);
INV_X1 g_I5801 (g1424, I5801);
INV_X1 g_g1923 (I5801, g1923);
INV_X1 g_g1924 (g174, g1924);
INV_X1 g_g1925 (g825, g1925);
INV_X1 g_g1926 (g874, g1926);
INV_X1 g_g1929 (g1224, g1929);
INV_X1 g_g1933 (g1247, g1933);
INV_X1 g_g1934 (g154, g1934);
INV_X1 g_g1935 (g1280, g1935);
INV_X1 g_g1938 (g1288, g1938);
INV_X1 g_I5812 (g1243, I5812);
INV_X1 g_g1941 (I5812, g1941);
INV_X1 g_g1942 (g828, g1942);
INV_X1 g_g1943 (g1025, g1943);
INV_X1 g_I5817 (g1081, I5817);
INV_X1 g_g1944 (I5817, g1944);
INV_X1 g_g1945 (g1081, g1945);
INV_X1 g_g1948 (g1250, g1948);
INV_X1 g_g1949 (g1292, g1949);
INV_X1 g_g1952 (g1333, g1952);
INV_X1 g_g1958 (g786, g1958);
INV_X1 g_g1959 (g1252, g1959);
INV_X1 g_g1960 (g1268, g1960);
INV_X1 g_g1961 (g1345, g1961);
INV_X1 g_g1967 (g1432, g1967);
INV_X1 g_I5831 (g1194, I5831);
INV_X1 g_g1970 (I5831, g1970);
INV_X1 g_g1974 (g803, g1974);
INV_X1 g_g1975 (g1253, g1975);
INV_X1 g_g1976 (g1269, g1976);
INV_X1 g_g1977 (g1357, g1977);
INV_X1 g_I5839 (g1198, I5839);
INV_X1 g_g1983 (I5839, g1983);
INV_X1 g_I5842 (g68, I5842);
INV_X1 g_g1987 (I5842, g1987);
INV_X1 g_g2006 (g806, g2006);
INV_X1 g_g2007 (g1223, g2007);
INV_X1 g_I5847 (g1360, I5847);
INV_X1 g_g2011 (I5847, g2011);
INV_X1 g_g2015 (g33, g2015);
INV_X1 g_I5852 (g1202, I5852);
INV_X1 g_g2016 (I5852, g2016);
INV_X1 g_I5855 (g71, I5855);
INV_X1 g_g2020 (I5855, g2020);
INV_X1 g_g2038 (g809, g2038);
INV_X1 g_g2039 (g1228, g2039);
INV_X1 g_I5861 (g1313, I5861);
INV_X1 g_g2044 (I5861, g2044);
INV_X1 g_I5865 (g1206, I5865);
INV_X1 g_g2052 (I5865, g2052);
INV_X1 g_I5868 (g74, I5868);
INV_X1 g_g2057 (I5868, g2057);
INV_X1 g_g2073 (g1254, g2073);
INV_X1 g_I5872 (g77, I5872);
INV_X1 g_g2074 (I5872, g2074);
INV_X1 g_g2091 (g819, g2091);
INV_X1 g_g2092 (g1225, g2092);
INV_X1 g_g2096 (g1226, g2096);
INV_X1 g_g2100 (g1227, g2100);
INV_X1 g_I5879 (g1267, I5879);
INV_X1 g_g2104 (I5879, g2104);
INV_X1 g_g2105 (g1444, g2105);
INV_X1 g_I5883 (g80, I5883);
INV_X1 g_g2106 (I5883, g2106);
INV_X1 g_g2128 (g1284, g2128);
INV_X1 g_g2131 (g1300, g2131);
INV_X1 g_g2134 (g1317, g2134);
INV_X1 g_I5889 (g83, I5889);
INV_X1 g_g2137 (I5889, g2137);
INV_X1 g_g2145 (g1296, g2145);
INV_X1 g_g2148 (g1304, g2148);
INV_X1 g_I5894 (g86, I5894);
INV_X1 g_g2149 (I5894, g2149);
INV_X1 g_I5897 (g173, I5897);
INV_X1 g_g2157 (I5897, g2157);
INV_X1 g_g2161 (g1454, g2161);
INV_X1 g_I5901 (g52, I5901);
INV_X1 g_g2162 (I5901, g2162);
INV_X1 g_g2170 (g1229, g2170);
INV_X1 g_g2174 (g1319, g2174);
INV_X1 g_g2177 (g1322, g2177);
INV_X1 g_g2180 (g1318, g2180);
INV_X1 g_I5908 (g196, I5908);
INV_X1 g_g2183 (I5908, g2183);
INV_X1 g_I5911 (g216, I5911);
INV_X1 g_g2184 (I5911, g2184);
INV_X1 g_I5914 (g1097, I5914);
INV_X1 g_g2185 (I5914, g2185);
INV_X1 g_g2202 (g1321, g2202);
INV_X1 g_g2205 (g13, g2205);
INV_X1 g_I5920 (g219, I5920);
INV_X1 g_g2207 (I5920, g2207);
INV_X1 g_I5923 (g252, I5923);
INV_X1 g_g2208 (I5923, g2208);
INV_X1 g_I5926 (g297, I5926);
INV_X1 g_g2209 (I5926, g2209);
INV_X1 g_g2210 (g1326, g2210);
INV_X1 g_g2215 (g1416, g2215);
INV_X1 g_I5933 (g1158, I5933);
INV_X1 g_g2216 (I5933, g2216);
INV_X1 g_I5936 (g222, I5936);
INV_X1 g_g2221 (I5936, g2221);
INV_X1 g_I5939 (g275, I5939);
INV_X1 g_g2222 (I5939, g2222);
INV_X1 g_I5942 (g300, I5942);
INV_X1 g_g2223 (I5942, g2223);
INV_X1 g_I5945 (g333, I5945);
INV_X1 g_g2224 (I5945, g2224);
INV_X1 g_I5948 (g378, I5948);
INV_X1 g_g2225 (I5948, g2225);
INV_X1 g_g2226 (g1320, g2226);
INV_X1 g_I5954 (g89, I5954);
INV_X1 g_g2231 (I5954, g2231);
INV_X1 g_I5957 (g110, I5957);
INV_X1 g_g2232 (I5957, g2232);
INV_X1 g_I5960 (g187, I5960);
INV_X1 g_g2233 (I5960, g2233);
INV_X1 g_I5963 (g225, I5963);
INV_X1 g_g2234 (I5963, g2234);
INV_X1 g_I5966 (g278, I5966);
INV_X1 g_g2235 (I5966, g2235);
INV_X1 g_I5969 (g303, I5969);
INV_X1 g_g2236 (I5969, g2236);
INV_X1 g_I5972 (g356, I5972);
INV_X1 g_g2237 (I5972, g2237);
INV_X1 g_I5975 (g381, I5975);
INV_X1 g_g2238 (I5975, g2238);
INV_X1 g_I5978 (g414, I5978);
INV_X1 g_g2239 (I5978, g2239);
INV_X1 g_I5981 (g459, I5981);
INV_X1 g_g2240 (I5981, g2240);
INV_X1 g_I5984 (g540, I5984);
INV_X1 g_g2241 (I5984, g2241);
INV_X1 g_g2242 (g985, g2242);
INV_X1 g_g2245 (g999, g2245);
INV_X1 g_I5989 (g1460, I5989);
INV_X1 g_g2246 (I5989, g2246);
INV_X1 g_g2253 (g1323, g2253);
INV_X1 g_g2256 (g1324, g2256);
INV_X1 g_g2259 (g1325, g2259);
INV_X1 g_g2263 (g1394, g2263);
INV_X1 g_I5997 (g114, I5997);
INV_X1 g_g2264 (I5997, g2264);
INV_X1 g_I6000 (g202, I6000);
INV_X1 g_g2265 (I6000, g2265);
INV_X1 g_I6003 (g228, I6003);
INV_X1 g_g2266 (I6003, g2266);
INV_X1 g_I6006 (g306, I6006);
INV_X1 g_g2267 (I6006, g2267);
INV_X1 g_I6009 (g359, I6009);
INV_X1 g_g2268 (I6009, g2268);
INV_X1 g_I6012 (g384, I6012);
INV_X1 g_g2269 (I6012, g2269);
INV_X1 g_I6015 (g437, I6015);
INV_X1 g_g2270 (I6015, g2270);
INV_X1 g_I6018 (g462, I6018);
INV_X1 g_g2271 (I6018, g2271);
INV_X1 g_I6021 (g495, I6021);
INV_X1 g_g2272 (I6021, g2272);
INV_X1 g_I6024 (g544, I6024);
INV_X1 g_g2273 (I6024, g2273);
INV_X1 g_g2274 (g782, g2274);
INV_X1 g_g2275 (g990, g2275);
INV_X1 g_I6029 (g1207, I6029);
INV_X1 g_g2276 (I6029, g2276);
INV_X1 g_g2282 (g1400, g2282);
INV_X1 g_I6033 (g3, I6033);
INV_X1 g_g2283 (I6033, g2283);
INV_X1 g_I6036 (g130, I6036);
INV_X1 g_g2284 (I6036, g2284);
INV_X1 g_I6039 (g207, I6039);
INV_X1 g_g2285 (I6039, g2285);
INV_X1 g_I6042 (g237, I6042);
INV_X1 g_g2286 (I6042, g2286);
INV_X1 g_I6045 (g309, I6045);
INV_X1 g_g2287 (I6045, g2287);
INV_X1 g_I6048 (g387, I6048);
INV_X1 g_g2288 (I6048, g2288);
INV_X1 g_I6051 (g440, I6051);
INV_X1 g_g2289 (I6051, g2289);
INV_X1 g_I6054 (g465, I6054);
INV_X1 g_g2290 (I6054, g2290);
INV_X1 g_I6057 (g518, I6057);
INV_X1 g_g2291 (I6057, g2291);
INV_X1 g_I6060 (g580, I6060);
INV_X1 g_g2292 (I6060, g2292);
INV_X1 g_g2293 (g888, g2293);
INV_X1 g_g2295 (g995, g2295);
INV_X1 g_I6072 (g1211, I6072);
INV_X1 g_g2298 (I6072, g2298);
INV_X1 g_I6075 (g2, I6075);
INV_X1 g_g2306 (I6075, g2306);
INV_X1 g_I6078 (g95, I6078);
INV_X1 g_g2307 (I6078, g2307);
INV_X1 g_I6081 (g118, I6081);
INV_X1 g_g2308 (I6081, g2308);
INV_X1 g_I6084 (g240, I6084);
INV_X1 g_g2309 (I6084, g2309);
INV_X1 g_I6087 (g318, I6087);
INV_X1 g_g2310 (I6087, g2310);
INV_X1 g_I6090 (g390, I6090);
INV_X1 g_g2311 (I6090, g2311);
INV_X1 g_I6093 (g468, I6093);
INV_X1 g_g2312 (I6093, g2312);
INV_X1 g_I6096 (g521, I6096);
INV_X1 g_g2313 (I6096, g2313);
INV_X1 g_I6099 (g584, I6099);
INV_X1 g_g2314 (I6099, g2314);
INV_X1 g_I6109 (g1214, I6109);
INV_X1 g_g2316 (I6109, g2316);
INV_X1 g_I6112 (g4, I6112);
INV_X1 g_g2323 (I6112, g2323);
INV_X1 g_I6115 (g134, I6115);
INV_X1 g_g2324 (I6115, g2324);
INV_X1 g_I6118 (g243, I6118);
INV_X1 g_g2325 (I6118, g2325);
INV_X1 g_I6121 (g321, I6121);
INV_X1 g_g2326 (I6121, g2326);
INV_X1 g_I6124 (g399, I6124);
INV_X1 g_g2327 (I6124, g2327);
INV_X1 g_I6127 (g471, I6127);
INV_X1 g_g2328 (I6127, g2328);
INV_X1 g_I6130 (g560, I6130);
INV_X1 g_g2329 (I6130, g2329);
INV_X1 g_g2331 (g933, g2331);
INV_X1 g_g2332 (g926, g2332);
INV_X1 g_I6143 (g1217, I6143);
INV_X1 g_g2334 (I6143, g2334);
INV_X1 g_g2340 (g1327, g2340);
INV_X1 g_g2343 (g1392, g2343);
INV_X1 g_I6148 (g5, I6148);
INV_X1 g_g2344 (I6148, g2344);
INV_X1 g_I6151 (g12, I6151);
INV_X1 g_g2345 (I6151, g2345);
INV_X1 g_I6154 (g122, I6154);
INV_X1 g_g2346 (I6154, g2346);
INV_X1 g_I6157 (g246, I6157);
INV_X1 g_g2347 (I6157, g2347);
INV_X1 g_I6160 (g324, I6160);
INV_X1 g_g2348 (I6160, g2348);
INV_X1 g_I6163 (g402, I6163);
INV_X1 g_g2349 (I6163, g2349);
INV_X1 g_I6166 (g480, I6166);
INV_X1 g_g2350 (I6166, g2350);
INV_X1 g_g2351 (g792, g2351);
INV_X1 g_g2353 (g871, g2353);
INV_X1 g_I6178 (g1220, I6178);
INV_X1 g_g2354 (I6178, g2354);
INV_X1 g_g2359 (g1397, g2359);
INV_X1 g_g2360 (g1435, g2360);
INV_X1 g_I6183 (g6, I6183);
INV_X1 g_g2361 (I6183, g2361);
INV_X1 g_I6186 (g138, I6186);
INV_X1 g_g2362 (I6186, g2362);
INV_X1 g_I6189 (g249, I6189);
INV_X1 g_g2363 (I6189, g2363);
INV_X1 g_I6192 (g327, I6192);
INV_X1 g_g2364 (I6192, g2364);
INV_X1 g_I6195 (g405, I6195);
INV_X1 g_g2365 (I6195, g2365);
INV_X1 g_I6198 (g483, I6198);
INV_X1 g_g2366 (I6198, g2366);
INV_X1 g_g2371 (g944, g2371);
INV_X1 g_I6214 (g7, I6214);
INV_X1 g_g2372 (I6214, g2372);
INV_X1 g_I6217 (g105, I6217);
INV_X1 g_g2373 (I6217, g2373);
INV_X1 g_I6220 (g126, I6220);
INV_X1 g_g2374 (I6220, g2374);
INV_X1 g_I6223 (g330, I6223);
INV_X1 g_g2375 (I6223, g2375);
INV_X1 g_I6226 (g408, I6226);
INV_X1 g_g2376 (I6226, g2376);
INV_X1 g_I6229 (g486, I6229);
INV_X1 g_g2377 (I6229, g2377);
INV_X1 g_I6239 (g8, I6239);
INV_X1 g_g2379 (I6239, g2379);
INV_X1 g_I6242 (g1554, I6242);
INV_X1 g_g2380 (I6242, g2380);
INV_X1 g_I6245 (g142, I6245);
INV_X1 g_g2381 (I6245, g2381);
INV_X1 g_I6248 (g411, I6248);
INV_X1 g_g2382 (I6248, g2382);
INV_X1 g_I6251 (g489, I6251);
INV_X1 g_g2383 (I6251, g2383);
INV_X1 g_I6254 (g536, I6254);
INV_X1 g_g2384 (I6254, g2384);
INV_X1 g_g2389 (g1230, g2389);
INV_X1 g_g2392 (g11, g2392);
INV_X1 g_I6267 (g100, I6267);
INV_X1 g_g2393 (I6267, g2393);
INV_X1 g_I6270 (g492, I6270);
INV_X1 g_g2394 (I6270, g2394);
INV_X1 g_g2396 (g1033, g2396);
INV_X1 g_g2397 (g1272, g2397);
INV_X1 g_g2401 (g22, g2401);
INV_X1 g_g2402 (g29, g2402);
INV_X1 g_g2403 (g1176, g2403);
INV_X1 g_g2404 (g1276, g2404);
INV_X1 g_I6286 (g1307, I6286);
INV_X1 g_g2407 (I6286, g2407);
INV_X1 g_g2424 (g1329, g2424);
INV_X1 g_g2452 (g23, g2452);
INV_X1 g_I6291 (g46, I6291);
INV_X1 g_g2453 (I6291, g2453);
INV_X1 g_I6294 (g1330, I6294);
INV_X1 g_g2454 (I6294, g2454);
INV_X1 g_g2457 (g24, g2457);
INV_X1 g_g2458 (g30, g2458);
INV_X1 g_I6299 (g47, I6299);
INV_X1 g_g2459 (I6299, g2459);
INV_X1 g_I6302 (g1313, I6302);
INV_X1 g_g2460 (I6302, g2460);
INV_X1 g_I6305 (g1333, I6305);
INV_X1 g_g2467 (I6305, g2467);
INV_X1 g_g2470 (g42, g2470);
INV_X1 g_I6309 (g1336, I6309);
INV_X1 g_g2471 (I6309, g2471);
INV_X1 g_g2477 (g25, g2477);
INV_X1 g_g2478 (g31, g2478);
INV_X1 g_g2479 (g32, g2479);
INV_X1 g_g2480 (g44, g2480);
INV_X1 g_I6317 (g1339, I6317);
INV_X1 g_g2481 (I6317, g2481);
INV_X1 g_g2484 (g45, g2484);
INV_X1 g_g2485 (g62, g2485);
INV_X1 g_g2486 (g959, g2486);
INV_X1 g_I6323 (g1342, I6323);
INV_X1 g_g2487 (I6323, g2487);
INV_X1 g_I6326 (g1443, I6326);
INV_X1 g_g2490 (I6326, g2490);
INV_X1 g_g2494 (g9, g2494);
INV_X1 g_g2495 (g26, g2495);
INV_X1 g_g2496 (g942, g2496);
INV_X1 g_g2497 (g945, g2497);
INV_X1 g_I6333 (g1345, I6333);
INV_X1 g_g2498 (I6333, g2498);
INV_X1 g_g2501 (g27, g2501);
INV_X1 g_I6337 (g1348, I6337);
INV_X1 g_g2502 (I6337, g2502);
INV_X1 g_g2505 (g28, g2505);
INV_X1 g_I6341 (g1351, I6341);
INV_X1 g_g2506 (I6341, g2506);
INV_X1 g_g2509 (g37, g2509);
INV_X1 g_g2510 (g58, g2510);
INV_X1 g_g2511 (g1328, g2511);
INV_X1 g_g2514 (g1330, g2514);
INV_X1 g_I6348 (g1354, I6348);
INV_X1 g_g2517 (I6348, g2517);
INV_X1 g_g2520 (g41, g2520);
INV_X1 g_g2522 (g1342, g2522);
INV_X1 g_I6354 (g1357, I6354);
INV_X1 g_g2525 (I6354, g2525);
INV_X1 g_g2528 (g1260, g2528);
INV_X1 g_I6358 (g13, I6358);
INV_X1 g_g2532 (I6358, g2532);
INV_X1 g_g2533 (g1336, g2533);
INV_X1 g_g2536 (g1354, g2536);
INV_X1 g_I6363 (g16, I6363);
INV_X1 g_g2539 (I6363, g2539);
INV_X1 g_g2540 (g1339, g2540);
INV_X1 g_g2543 (g1348, g2543);
INV_X1 g_I6368 (g20, I6368);
INV_X1 g_g2546 (I6368, g2546);
INV_X1 g_I6371 (g33, I6371);
INV_X1 g_g2547 (I6371, g2547);
INV_X1 g_g2548 (g1351, g2548);
INV_X1 g_g2551 (g1360, g2551);
INV_X1 g_I6376 (g38, I6376);
INV_X1 g_g2554 (I6376, g2554);
INV_X1 g_g2555 (g936, g2555);
INV_X1 g_g2556 (g1190, g2556);
INV_X1 g_g2557 (g940, g2557);
INV_X1 g_g2561 (g1555, g2561);
INV_X1 g_g2562 (g1652, g2562);
INV_X1 g_g2573 (g1649, g2573);
INV_X1 g_g2584 (g1646, g2584);
INV_X1 g_g2595 (g1643, g2595);
INV_X1 g_g2605 (g1639, g2605);
INV_X1 g_g2614 (g1562, g2614);
INV_X1 g_g2615 (g1563, g2615);
INV_X1 g_g2616 (g1564, g2616);
INV_X1 g_g2617 (g1565, g2617);
INV_X1 g_g2618 (g1566, g2618);
INV_X1 g_g2621 (g1567, g2621);
INV_X1 g_g2622 (g1568, g2622);
INV_X1 g_g2623 (g1585, g2623);
INV_X1 g_g2624 (g1569, g2624);
INV_X1 g_g2625 (g1570, g2625);
INV_X1 g_g2626 (g1571, g2626);
INV_X1 g_g2627 (g1572, g2627);
INV_X1 g_g2628 (g1573, g2628);
INV_X1 g_g2629 (g1574, g2629);
INV_X1 g_g2630 (g1575, g2630);
INV_X1 g_g2631 (g1586, g2631);
INV_X1 g_g2632 (g1576, g2632);
INV_X1 g_g2633 (g1577, g2633);
INV_X1 g_g2634 (g1578, g2634);
INV_X1 g_g2635 (g1579, g2635);
INV_X1 g_g2636 (g1580, g2636);
INV_X1 g_g2637 (g1581, g2637);
INV_X1 g_g2638 (g1582, g2638);
INV_X1 g_g2639 (g1583, g2639);
INV_X1 g_g2640 (g1584, g2640);
INV_X1 g_g2641 (g1587, g2641);
INV_X1 g_g2642 (g1588, g2642);
INV_X1 g_g2643 (g1589, g2643);
INV_X1 g_I6416 (g1794, I6416);
INV_X1 g_g2644 (I6416, g2644);
INV_X1 g_I6419 (g1799, I6419);
INV_X1 g_g2645 (I6419, g2645);
INV_X1 g_I6422 (g1805, I6422);
INV_X1 g_g2646 (I6422, g2646);
INV_X1 g_I6425 (g1811, I6425);
INV_X1 g_g2647 (I6425, g2647);
INV_X1 g_I6428 (g1818, I6428);
INV_X1 g_g2648 (I6428, g2648);
INV_X1 g_I6431 (g1825, I6431);
INV_X1 g_g2649 (I6431, g2649);
INV_X1 g_I6434 (g1830, I6434);
INV_X1 g_g2650 (I6434, g2650);
INV_X1 g_I6437 (g1784, I6437);
INV_X1 g_g2651 (I6437, g2651);
INV_X1 g_I6440 (g1806, I6440);
INV_X1 g_g2652 (I6440, g2652);
INV_X1 g_I6443 (g1774, I6443);
INV_X1 g_g2653 (I6443, g2653);
INV_X1 g_I6446 (g1812, I6446);
INV_X1 g_g2654 (I6446, g2654);
INV_X1 g_g2655 (g1611, g2655);
INV_X1 g_g2659 (g1655, g2659);
INV_X1 g_I6451 (g1895, I6451);
INV_X1 g_g2660 (I6451, g2660);
INV_X1 g_I6454 (g1868, I6454);
INV_X1 g_g2661 (I6454, g2661);
INV_X1 g_I6457 (g1886, I6457);
INV_X1 g_g2662 (I6457, g2662);
INV_X1 g_I6460 (g2104, I6460);
INV_X1 g_g2663 (I6460, g2663);
INV_X1 g_I6463 (g1769, I6463);
INV_X1 g_g2664 (I6463, g2664);
INV_X1 g_g2665 (g1661, g2665);
INV_X1 g_g2668 (g1662, g2668);
INV_X1 g_I6468 (g1917, I6468);
INV_X1 g_g2671 (I6468, g2671);
INV_X1 g_I6471 (g1923, I6471);
INV_X1 g_g2672 (I6471, g2672);
INV_X1 g_I6474 (g1941, I6474);
INV_X1 g_g2673 (I6474, g2673);
INV_X1 g_g2674 (g1675, g2674);
INV_X1 g_g2677 (g1664, g2677);
INV_X1 g_g2680 (g1665, g2680);
INV_X1 g_g2683 (g1666, g2683);
INV_X1 g_g2686 (g1667, g2686);
INV_X1 g_g2689 (g1670, g2689);
INV_X1 g_g2692 (g1671, g2692);
INV_X1 g_g2695 (g1672, g2695);
INV_X1 g_g2698 (g1673, g2698);
INV_X1 g_g2699 (g1674, g2699);
INV_X1 g_g2700 (g1744, g2700);
INV_X1 g_g2703 (g1809, g2703);
INV_X1 g_g2706 (g1821, g2706);
INV_X1 g_g2709 (g1747, g2709);
INV_X1 g_g2712 (g2039, g2712);
INV_X1 g_g2721 (g1803, g2721);
INV_X1 g_g2724 (g1814, g2724);
INV_X1 g_g2727 (g2424, g2727);
INV_X1 g_g2728 (g2256, g2728);
INV_X1 g_g2734 (g2170, g2734);
INV_X1 g_g2743 (g1808, g2743);
INV_X1 g_g2746 (g2259, g2746);
INV_X1 g_g2752 (g2389, g2752);
INV_X1 g_g2761 (g1820, g2761);
INV_X1 g_g2764 (g1802, g2764);
INV_X1 g_I6509 (g1684, I6509);
INV_X1 g_g2767 (I6509, g2767);
INV_X1 g_g2769 (g2424, g2769);
INV_X1 g_g2770 (g2210, g2770);
INV_X1 g_g2774 (g1813, g2774);
INV_X1 g_g2777 (g1797, g2777);
INV_X1 g_I6517 (g1687, I6517);
INV_X1 g_g2780 (I6517, g2780);
INV_X1 g_g2782 (g1616, g2782);
INV_X1 g_g2784 (g2340, g2784);
INV_X1 g_g2787 (g1807, g2787);
INV_X1 g_g2790 (g1793, g2790);
INV_X1 g_I6532 (g1694, I6532);
INV_X1 g_g2793 (I6532, g2793);
INV_X1 g_g2794 (g2185, g2794);
INV_X1 g_g2795 (g1801, g2795);
INV_X1 g_g2798 (g1787, g2798);
INV_X1 g_g2804 (g1796, g2804);
INV_X1 g_g2807 (g1782, g2807);
INV_X1 g_g2810 (g1922, g2810);
INV_X1 g_g2816 (g1685, g2816);
INV_X1 g_g2817 (g1849, g2817);
INV_X1 g_g2818 (g1792, g2818);
INV_X1 g_g2821 (g1786, g2821);
INV_X1 g_g2824 (g1688, g2824);
INV_X1 g_I6553 (g2246, I6553);
INV_X1 g_g2825 (I6553, g2825);
INV_X1 g_g2826 (g2183, g2826);
INV_X1 g_g2828 (g1980, g2828);
INV_X1 g_g2829 (g1785, g2829);
INV_X1 g_g2832 (g2184, g2832);
INV_X1 g_I6561 (g1715, I6561);
INV_X1 g_g2833 (I6561, g2833);
INV_X1 g_I6564 (g2073, I6564);
INV_X1 g_g2834 (I6564, g2834);
INV_X1 g_g2837 (g1780, g2837);
INV_X1 g_g2840 (g2207, g2840);
INV_X1 g_g2841 (g2208, g2841);
INV_X1 g_g2842 (g2209, g2842);
INV_X1 g_I6571 (g1711, I6571);
INV_X1 g_g2843 (I6571, g2843);
INV_X1 g_I6574 (g576, I6574);
INV_X1 g_g2844 (I6574, g2844);
INV_X1 g_I6578 (g1603, I6578);
INV_X1 g_g2862 (I6578, g2862);
INV_X1 g_g2863 (g1778, g2863);
INV_X1 g_g2866 (g2221, g2866);
INV_X1 g_g2867 (g2222, g2867);
INV_X1 g_g2868 (g2223, g2868);
INV_X1 g_g2869 (g2224, g2869);
INV_X1 g_g2870 (g2225, g2870);
INV_X1 g_I6587 (g1708, I6587);
INV_X1 g_g2871 (I6587, g2871);
INV_X1 g_I6590 (g2467, I6590);
INV_X1 g_g2872 (I6590, g2872);
INV_X1 g_g2873 (g1779, g2873);
INV_X1 g_g2876 (g2231, g2876);
INV_X1 g_g2877 (g2232, g2877);
INV_X1 g_g2878 (g2233, g2878);
INV_X1 g_I6597 (g1970, I6597);
INV_X1 g_g2879 (I6597, g2879);
INV_X1 g_g2880 (g2234, g2880);
INV_X1 g_g2881 (g2235, g2881);
INV_X1 g_g2882 (g2236, g2882);
INV_X1 g_g2883 (g2237, g2883);
INV_X1 g_g2884 (g2238, g2884);
INV_X1 g_g2885 (g2239, g2885);
INV_X1 g_g2886 (g2240, g2886);
INV_X1 g_g2887 (g2241, g2887);
INV_X1 g_I6608 (g1612, I6608);
INV_X1 g_g2888 (I6608, g2888);
INV_X1 g_g2890 (g2264, g2890);
INV_X1 g_g2891 (g2265, g2891);
INV_X1 g_g2892 (g2266, g2892);
INV_X1 g_I6615 (g1983, I6615);
INV_X1 g_g2893 (I6615, g2893);
INV_X1 g_g2894 (g2267, g2894);
INV_X1 g_g2895 (g2268, g2895);
INV_X1 g_g2896 (g2269, g2896);
INV_X1 g_g2897 (g2270, g2897);
INV_X1 g_g2898 (g2271, g2898);
INV_X1 g_g2899 (g2272, g2899);
INV_X1 g_g2900 (g2273, g2900);
INV_X1 g_g2901 (g2284, g2901);
INV_X1 g_g2902 (g2285, g2902);
INV_X1 g_g2903 (g2286, g2903);
INV_X1 g_g2904 (g2287, g2904);
INV_X1 g_I6629 (g2052, I6629);
INV_X1 g_g2905 (I6629, g2905);
INV_X1 g_g2906 (g2288, g2906);
INV_X1 g_g2907 (g2289, g2907);
INV_X1 g_g2908 (g2290, g2908);
INV_X1 g_g2909 (g2291, g2909);
INV_X1 g_I6636 (g1704, I6636);
INV_X1 g_g2910 (I6636, g2910);
INV_X1 g_g2911 (g2292, g2911);
INV_X1 g_g2913 (g2307, g2913);
INV_X1 g_g2914 (g2308, g2914);
INV_X1 g_I6643 (g1970, I6643);
INV_X1 g_g2915 (I6643, g2915);
INV_X1 g_I6646 (g2246, I6646);
INV_X1 g_g2916 (I6646, g2916);
INV_X1 g_g2917 (g2309, g2917);
INV_X1 g_g2918 (g2310, g2918);
INV_X1 g_g2919 (g2311, g2919);
INV_X1 g_I6652 (g2016, I6652);
INV_X1 g_g2920 (I6652, g2920);
INV_X1 g_g2921 (g2312, g2921);
INV_X1 g_g2922 (g2313, g2922);
INV_X1 g_I6657 (g1701, I6657);
INV_X1 g_g2923 (I6657, g2923);
INV_X1 g_g2924 (g2314, g2924);
INV_X1 g_g2925 (g2324, g2925);
INV_X1 g_g2926 (g2325, g2926);
INV_X1 g_I6663 (g2246, I6663);
INV_X1 g_g2927 (I6663, g2927);
INV_X1 g_g2928 (g2326, g2928);
INV_X1 g_g2929 (g2327, g2929);
INV_X1 g_g2930 (g2328, g2930);
INV_X1 g_I6669 (g1698, I6669);
INV_X1 g_g2931 (I6669, g2931);
INV_X1 g_g2932 (g2329, g2932);
INV_X1 g_I6673 (g2246, I6673);
INV_X1 g_g2933 (I6673, g2933);
INV_X1 g_I6676 (g1603, I6676);
INV_X1 g_g2934 (I6676, g2934);
INV_X1 g_I6680 (g1558, I6680);
INV_X1 g_g2936 (I6680, g2936);
INV_X1 g_g2937 (g2346, g2937);
INV_X1 g_g2938 (g2347, g2938);
INV_X1 g_g2939 (g2348, g2939);
INV_X1 g_I6686 (g2246, I6686);
INV_X1 g_g2940 (I6686, g2940);
INV_X1 g_g2941 (g2349, g2941);
INV_X1 g_g2942 (g2350, g2942);
INV_X1 g_g2943 (g2362, g2943);
INV_X1 g_g2944 (g2363, g2944);
INV_X1 g_g2945 (g2364, g2945);
INV_X1 g_g2946 (g2365, g2946);
INV_X1 g_I6695 (g2246, I6695);
INV_X1 g_g2947 (I6695, g2947);
INV_X1 g_g2948 (g2366, g2948);
INV_X1 g_g2953 (g2373, g2953);
INV_X1 g_g2954 (g2374, g2954);
INV_X1 g_I6703 (g1983, I6703);
INV_X1 g_g2955 (I6703, g2955);
INV_X1 g_g2956 (g2375, g2956);
INV_X1 g_g2957 (g2376, g2957);
INV_X1 g_g2958 (g2377, g2958);
INV_X1 g_g2959 (g1926, g2959);
INV_X1 g_g2960 (g2381, g2960);
INV_X1 g_I6711 (g1726, I6711);
INV_X1 g_g2961 (I6711, g2961);
INV_X1 g_g2962 (g2382, g2962);
INV_X1 g_g2963 (g2383, g2963);
INV_X1 g_I6716 (g1721, I6716);
INV_X1 g_g2964 (I6716, g2964);
INV_X1 g_g2965 (g2384, g2965);
INV_X1 g_g2966 (g1856, g2966);
INV_X1 g_g2969 (g2393, g2969);
INV_X1 g_g2970 (g2394, g2970);
INV_X1 g_I6723 (g2052, I6723);
INV_X1 g_g2971 (I6723, g2971);
INV_X1 g_g2973 (g1854, g2973);
INV_X1 g_I6728 (g1959, I6728);
INV_X1 g_g2976 (I6728, g2976);
INV_X1 g_g2982 (g1848, g2982);
INV_X1 g_I6733 (g1718, I6733);
INV_X1 g_g2985 (I6733, g2985);
INV_X1 g_g2989 (g1843, g2989);
INV_X1 g_g2992 (g1833, g2992);
INV_X1 g_g2996 (g1828, g2996);
INV_X1 g_g2999 (g1823, g2999);
INV_X1 g_g3008 (g1816, g3008);
INV_X1 g_I6764 (g1955, I6764);
INV_X1 g_g3013 (I6764, g3013);
INV_X1 g_I6767 (g1933, I6767);
INV_X1 g_g3014 (I6767, g3014);
INV_X1 g_I6770 (g1590, I6770);
INV_X1 g_g3018 (I6770, g3018);
INV_X1 g_g3019 (g2007, g3019);
INV_X1 g_g3029 (g1929, g3029);
INV_X1 g_g3038 (g2092, g3038);
INV_X1 g_g3047 (g1736, g3047);
INV_X1 g_I6784 (g2052, I6784);
INV_X1 g_g3048 (I6784, g3048);
INV_X1 g_I6788 (g1681, I6788);
INV_X1 g_g3050 (I6788, g3050);
INV_X1 g_I6791 (g1967, I6791);
INV_X1 g_g3051 (I6791, g3051);
INV_X1 g_g3052 (g2096, g3052);
INV_X1 g_I6795 (g1683, I6795);
INV_X1 g_g3061 (I6795, g3061);
INV_X1 g_g3062 (g2100, g3062);
INV_X1 g_g3071 (g1948, g3071);
INV_X1 g_I6800 (g2016, I6800);
INV_X1 g_g3074 (I6800, g3074);
INV_X1 g_g3075 (g2216, g3075);
INV_X1 g_g3076 (g1831, g3076);
INV_X1 g_I6805 (g1603, I6805);
INV_X1 g_g3077 (I6805, g3077);
INV_X1 g_g3078 (g1603, g3078);
INV_X1 g_g3079 (g1603, g3079);
INV_X1 g_g3080 (g1679, g3080);
INV_X1 g_g3082 (g1680, g3082);
INV_X1 g_I6820 (g1707, I6820);
INV_X1 g_g3084 (I6820, g3084);
INV_X1 g_g3085 (g1945, g3085);
INV_X1 g_g3086 (g1852, g3086);
INV_X1 g_g3091 (g1603, g3091);
INV_X1 g_I6826 (g2185, I6826);
INV_X1 g_g3092 (I6826, g3092);
INV_X1 g_g3093 (g1686, g3093);
INV_X1 g_I6831 (g2185, I6831);
INV_X1 g_g3095 (I6831, g3095);
INV_X1 g_I6834 (g287, I6834);
INV_X1 g_g3096 (I6834, g3096);
INV_X1 g_g3124 (g1857, g3124);
INV_X1 g_I6839 (g2185, I6839);
INV_X1 g_g3128 (I6839, g3128);
INV_X1 g_I6849 (g368, I6849);
INV_X1 g_g3130 (I6849, g3130);
INV_X1 g_I6853 (g2185, I6853);
INV_X1 g_g3158 (I6853, g3158);
INV_X1 g_I6856 (g449, I6856);
INV_X1 g_g3159 (I6856, g3159);
INV_X1 g_I6860 (g2185, I6860);
INV_X1 g_g3187 (I6860, g3187);
INV_X1 g_I6864 (g2528, I6864);
INV_X1 g_g3189 (I6864, g3189);
INV_X1 g_I6868 (g530, I6868);
INV_X1 g_g3191 (I6868, g3191);
INV_X1 g_I6872 (g2185, I6872);
INV_X1 g_g3219 (I6872, g3219);
INV_X1 g_g3220 (g1889, g3220);
INV_X1 g_I6887 (g2528, I6887);
INV_X1 g_g3230 (I6887, g3230);
INV_X1 g_I6894 (g1863, I6894);
INV_X1 g_g3238 (I6894, g3238);
INV_X1 g_I6900 (g1866, I6900);
INV_X1 g_g3264 (I6900, g3264);
INV_X1 g_g3285 (g1689, g3285);
INV_X1 g_I6911 (g1869, I6911);
INV_X1 g_g3287 (I6911, g3287);
INV_X1 g_I6930 (g1876, I6930);
INV_X1 g_g3316 (I6930, g3316);
INV_X1 g_g3338 (g1901, g3338);
INV_X1 g_g3340 (g2474, g3340);
INV_X1 g_I6936 (g1878, I6936);
INV_X1 g_g3341 (I6936, g3341);
INV_X1 g_I6946 (g1887, I6946);
INV_X1 g_g3359 (I6946, g3359);
INV_X1 g_I6949 (g2148, I6949);
INV_X1 g_g3390 (I6949, g3390);
INV_X1 g_I6952 (g1896, I6952);
INV_X1 g_g3398 (I6952, g3398);
INV_X1 g_I6956 (g1907, I6956);
INV_X1 g_g3430 (I6956, g3430);
INV_X1 g_I6959 (g1558, I6959);
INV_X1 g_g3461 (I6959, g3461);
INV_X1 g_g3462 (g1743, g3462);
INV_X1 g_I6963 (g1558, I6963);
INV_X1 g_g3465 (I6963, g3465);
INV_X1 g_g3485 (g1737, g3485);
INV_X1 g_g3488 (g1727, g3488);
INV_X1 g_g3491 (g1800, g3491);
INV_X1 g_I6970 (g1872, I6970);
INV_X1 g_g3492 (I6970, g3492);
INV_X1 g_g3495 (g1616, g3495);
INV_X1 g_I6974 (g2528, I6974);
INV_X1 g_g3496 (I6974, g3496);
INV_X1 g_g3497 (g2185, g3497);
INV_X1 g_g3498 (g1616, g3498);
INV_X1 g_g3499 (g2185, g3499);
INV_X1 g_g3500 (g1616, g3500);
INV_X1 g_g3501 (g2185, g3501);
INV_X1 g_g3502 (g1616, g3502);
INV_X1 g_g3503 (g2407, g3503);
INV_X1 g_g3506 (g1781, g3506);
INV_X1 g_g3510 (g2185, g3510);
INV_X1 g_g3511 (g1616, g3511);
INV_X1 g_g3512 (g1616, g3512);
INV_X1 g_g3513 (g2407, g3513);
INV_X1 g_g3514 (g2424, g3514);
INV_X1 g_g3517 (g2283, g3517);
INV_X1 g_g3519 (g2185, g3519);
INV_X1 g_g3520 (g1616, g3520);
INV_X1 g_g3521 (g2185, g3521);
INV_X1 g_g3522 (g2407, g3522);
INV_X1 g_g3523 (g2407, g3523);
INV_X1 g_g3524 (g2306, g3524);
INV_X1 g_g3526 (g2185, g3526);
INV_X1 g_g3527 (g1616, g3527);
INV_X1 g_g3529 (g2323, g3529);
INV_X1 g_g3530 (g2185, g3530);
INV_X1 g_g3531 (g1616, g3531);
INV_X1 g_g3532 (g2407, g3532);
INV_X1 g_g3533 (g2397, g3533);
INV_X1 g_g3539 (g2424, g3539);
INV_X1 g_g3540 (g2424, g3540);
INV_X1 g_g3542 (g1777, g3542);
INV_X1 g_g3545 (g2344, g3545);
INV_X1 g_I7029 (g2392, I7029);
INV_X1 g_g3546 (I7029, g3546);
INV_X1 g_g3547 (g2345, g3547);
INV_X1 g_g3548 (g2185, g3548);
INV_X1 g_g3549 (g2404, g3549);
INV_X1 g_I7036 (g2454, I7036);
INV_X1 g_g3556 (I7036, g3556);
INV_X1 g_g3557 (g1773, g3557);
INV_X1 g_g3560 (g2361, g3560);
INV_X1 g_I7041 (g2401, I7041);
INV_X1 g_g3561 (I7041, g3561);
INV_X1 g_I7044 (g2402, I7044);
INV_X1 g_g3562 (I7044, g3562);
INV_X1 g_g3563 (g2007, g3563);
INV_X1 g_g3567 (g2407, g3567);
INV_X1 g_g3568 (g1935, g3568);
INV_X1 g_g3573 (g2424, g3573);
INV_X1 g_g3574 (g1771, g3574);
INV_X1 g_g3577 (g2372, g3577);
INV_X1 g_I7053 (g2452, I7053);
INV_X1 g_g3578 (I7053, g3578);
INV_X1 g_g3579 (g1929, g3579);
INV_X1 g_g3582 (g2407, g3582);
INV_X1 g_g3583 (g2128, g3583);
INV_X1 g_g3587 (g1964, g3587);
INV_X1 g_g3588 (g2379, g3588);
INV_X1 g_I7061 (g2457, I7061);
INV_X1 g_g3589 (I7061, g3589);
INV_X1 g_I7064 (g2458, I7064);
INV_X1 g_g3590 (I7064, g3590);
INV_X1 g_g3591 (g1789, g3591);
INV_X1 g_g3603 (g2092, g3603);
INV_X1 g_g3604 (g2407, g3604);
INV_X1 g_g3605 (g1938, g3605);
INV_X1 g_g3610 (g2424, g3610);
INV_X1 g_I7079 (g2532, I7079);
INV_X1 g_g3611 (I7079, g3611);
INV_X1 g_I7082 (g2470, I7082);
INV_X1 g_g3612 (I7082, g3612);
INV_X1 g_g3617 (g1655, g3617);
INV_X1 g_g3629 (g2424, g3629);
INV_X1 g_I7095 (g2539, I7095);
INV_X1 g_g3630 (I7095, g3630);
INV_X1 g_I7098 (g2477, I7098);
INV_X1 g_g3631 (I7098, g3631);
INV_X1 g_I7101 (g2478, I7101);
INV_X1 g_g3632 (I7101, g3632);
INV_X1 g_I7104 (g2479, I7104);
INV_X1 g_g3633 (I7104, g3633);
INV_X1 g_I7107 (g2480, I7107);
INV_X1 g_g3634 (I7107, g3634);
INV_X1 g_g3635 (g1949, g3635);
INV_X1 g_g3639 (g2424, g3639);
INV_X1 g_I7112 (g2546, I7112);
INV_X1 g_g3640 (I7112, g3640);
INV_X1 g_I7115 (g2547, I7115);
INV_X1 g_g3641 (I7115, g3641);
INV_X1 g_I7118 (g2484, I7118);
INV_X1 g_g3642 (I7118, g3642);
INV_X1 g_g3643 (g2453, g3643);
INV_X1 g_g3644 (g2131, g3644);
INV_X1 g_g3647 (g2424, g3647);
INV_X1 g_g3648 (g2424, g3648);
INV_X1 g_g3649 (g2424, g3649);
INV_X1 g_I7126 (g2494, I7126);
INV_X1 g_g3650 (I7126, g3650);
INV_X1 g_I7129 (g2495, I7129);
INV_X1 g_g3651 (I7129, g3651);
INV_X1 g_I7132 (g2554, I7132);
INV_X1 g_g3652 (I7132, g3652);
INV_X1 g_g3653 (g2459, g3653);
INV_X1 g_g3654 (g2521, g3654);
INV_X1 g_g3655 (g1844, g3655);
INV_X1 g_I7145 (g2501, I7145);
INV_X1 g_g3657 (I7145, g3657);
INV_X1 g_g3659 (g2293, g3659);
INV_X1 g_g3666 (g2134, g3666);
INV_X1 g_I7164 (g2157, I7164);
INV_X1 g_g3674 (I7164, g3674);
INV_X1 g_I7167 (g2505, I7167);
INV_X1 g_g3675 (I7167, g3675);
INV_X1 g_g3676 (g2380, g3676);
INV_X1 g_g3677 (g2485, g3677);
INV_X1 g_g3684 (g2180, g3684);
INV_X1 g_I7195 (g1795, I7195);
INV_X1 g_g3691 (I7195, g3691);
INV_X1 g_I7198 (g2509, I7198);
INV_X1 g_g3692 (I7198, g3692);
INV_X1 g_g3693 (g2424, g3693);
INV_X1 g_g3694 (g2174, g3694);
INV_X1 g_g3700 (g2514, g3700);
INV_X1 g_I7204 (g2520, I7204);
INV_X1 g_g3705 (I7204, g3705);
INV_X1 g_g3707 (g2226, g3707);
INV_X1 g_g3712 (g1952, g3712);
INV_X1 g_g3716 (g2522, g3716);
INV_X1 g_I7211 (g1742, I7211);
INV_X1 g_g3721 (I7211, g3721);
INV_X1 g_g3723 (g2096, g3723);
INV_X1 g_g3728 (g2202, g3728);
INV_X1 g_g3732 (g2533, g3732);
INV_X1 g_g3735 (g1961, g3735);
INV_X1 g_g3739 (g2536, g3739);
INV_X1 g_g3743 (g1776, g3743);
INV_X1 g_g3746 (g2100, g3746);
INV_X1 g_g3750 (g2177, g3750);
INV_X1 g_g3753 (g2540, g3753);
INV_X1 g_g3754 (g2543, g3754);
INV_X1 g_g3757 (g1977, g3757);
INV_X1 g_g3761 (g1772, g3761);
INV_X1 g_g3764 (g2039, g3764);
INV_X1 g_g3768 (g2253, g3768);
INV_X1 g_g3769 (g2548, g3769);
INV_X1 g_g3770 (g2551, g3770);
INV_X1 g_g3771 (g1853, g3771);
INV_X1 g_g3774 (g1770, g3774);
INV_X1 g_g3777 (g2170, g3777);
INV_X1 g_g3778 (g2145, g3778);
INV_X1 g_g3779 (g2511, g3779);
INV_X1 g_g3780 (g1847, g3780);
INV_X1 g_I7255 (g1955, I7255);
INV_X1 g_g3783 (I7255, g3783);
INV_X1 g_g3784 (g1768, g3784);
INV_X1 g_g3787 (g1842, g3787);
INV_X1 g_g3798 (g1757, g3798);
INV_X1 g_I7262 (g2514, I7262);
INV_X1 g_g3801 (I7262, g3801);
INV_X1 g_g3802 (g1832, g3802);
INV_X1 g_g3805 (g1752, g3805);
INV_X1 g_g3808 (g1827, g3808);
INV_X1 g_g3812 (g1750, g3812);
INV_X1 g_g3815 (g1822, g3815);
INV_X1 g_g3819 (g1748, g3819);
INV_X1 g_g3822 (g1815, g3822);
INV_X1 g_g3825 (g1826, g3825);
INV_X1 g_I7287 (g2561, I7287);
INV_X1 g_g3828 (I7287, g3828);
INV_X1 g_I7290 (g2936, I7290);
INV_X1 g_g3829 (I7290, g3829);
INV_X1 g_I7293 (g2955, I7293);
INV_X1 g_g3830 (I7293, g3830);
INV_X1 g_I7296 (g2915, I7296);
INV_X1 g_g3831 (I7296, g3831);
INV_X1 g_I7299 (g2961, I7299);
INV_X1 g_g3832 (I7299, g3832);
INV_X1 g_I7302 (g2825, I7302);
INV_X1 g_g3833 (I7302, g3833);
INV_X1 g_I7305 (g3048, I7305);
INV_X1 g_g3834 (I7305, g3834);
INV_X1 g_I7308 (g3074, I7308);
INV_X1 g_g3835 (I7308, g3835);
INV_X1 g_I7311 (g2879, I7311);
INV_X1 g_g3836 (I7311, g3836);
INV_X1 g_I7314 (g2916, I7314);
INV_X1 g_g3837 (I7314, g3837);
INV_X1 g_I7317 (g2893, I7317);
INV_X1 g_g3838 (I7317, g3838);
INV_X1 g_I7320 (g2927, I7320);
INV_X1 g_g3839 (I7320, g3839);
INV_X1 g_I7323 (g2905, I7323);
INV_X1 g_g3840 (I7323, g3840);
INV_X1 g_I7326 (g2940, I7326);
INV_X1 g_g3841 (I7326, g3841);
INV_X1 g_I7329 (g2920, I7329);
INV_X1 g_g3842 (I7329, g3842);
INV_X1 g_I7332 (g2947, I7332);
INV_X1 g_g3843 (I7332, g3843);
INV_X1 g_I7335 (g2910, I7335);
INV_X1 g_g3844 (I7335, g3844);
INV_X1 g_I7338 (g2923, I7338);
INV_X1 g_g3845 (I7338, g3845);
INV_X1 g_I7341 (g2931, I7341);
INV_X1 g_g3846 (I7341, g3846);
INV_X1 g_I7344 (g2964, I7344);
INV_X1 g_g3847 (I7344, g3847);
INV_X1 g_I7347 (g2985, I7347);
INV_X1 g_g3848 (I7347, g3848);
INV_X1 g_I7350 (g2971, I7350);
INV_X1 g_g3849 (I7350, g3849);
INV_X1 g_I7353 (g2833, I7353);
INV_X1 g_g3850 (I7353, g3850);
INV_X1 g_I7356 (g2843, I7356);
INV_X1 g_g3851 (I7356, g3851);
INV_X1 g_I7359 (g2871, I7359);
INV_X1 g_g3852 (I7359, g3852);
INV_X1 g_I7362 (g2933, I7362);
INV_X1 g_g3853 (I7362, g3853);
INV_X1 g_I7365 (g3061, I7365);
INV_X1 g_g3854 (I7365, g3854);
INV_X1 g_I7368 (g3018, I7368);
INV_X1 g_g3855 (I7368, g3855);
INV_X1 g_I7371 (g3050, I7371);
INV_X1 g_g3856 (I7371, g3856);
INV_X1 g_I7374 (g3084, I7374);
INV_X1 g_g3857 (I7374, g3857);
INV_X1 g_I7377 (g3189, I7377);
INV_X1 g_g3858 (I7377, g3858);
INV_X1 g_I7380 (g3461, I7380);
INV_X1 g_g3859 (I7380, g3859);
INV_X1 g_I7383 (g3465, I7383);
INV_X1 g_g3860 (I7383, g3860);
INV_X1 g_I7386 (g3013, I7386);
INV_X1 g_g3861 (I7386, g3861);
INV_X1 g_I7389 (g3496, I7389);
INV_X1 g_g3862 (I7389, g3862);
INV_X1 g_I7392 (g3230, I7392);
INV_X1 g_g3863 (I7392, g3863);
INV_X1 g_g3864 (g2943, g3864);
INV_X1 g_g3865 (g2944, g3865);
INV_X1 g_g3866 (g2945, g3866);
INV_X1 g_g3867 (g2946, g3867);
INV_X1 g_g3868 (g2948, g3868);
INV_X1 g_I7400 (g3075, I7400);
INV_X1 g_g3869 (I7400, g3869);
INV_X1 g_g3870 (g3466, g3870);
INV_X1 g_g3871 (g2953, g3871);
INV_X1 g_g3872 (g2954, g3872);
INV_X1 g_g3873 (g2956, g3873);
INV_X1 g_g3874 (g2957, g3874);
INV_X1 g_g3875 (g2958, g3875);
INV_X1 g_g3876 (g3466, g3876);
INV_X1 g_g3877 (g2960, g3877);
INV_X1 g_g3878 (g2962, g3878);
INV_X1 g_g3879 (g2963, g3879);
INV_X1 g_g3880 (g2965, g3880);
INV_X1 g_g3881 (g2969, g3881);
INV_X1 g_g3882 (g2970, g3882);
INV_X1 g_I7417 (g3659, I7417);
INV_X1 g_g3884 (I7417, g3884);
INV_X1 g_g3888 (g3097, g3888);
INV_X1 g_g3891 (g3097, g3891);
INV_X1 g_g3892 (g3131, g3892);
INV_X1 g_I7473 (g3546, I7473);
INV_X1 g_g3896 (I7473, g3896);
INV_X1 g_g3897 (g3131, g3897);
INV_X1 g_g3898 (g3160, g3898);
INV_X1 g_I7492 (g3561, I7492);
INV_X1 g_g3901 (I7492, g3901);
INV_X1 g_I7495 (g3562, I7495);
INV_X1 g_g3902 (I7495, g3902);
INV_X1 g_I7498 (g2752, I7498);
INV_X1 g_g3903 (I7498, g3903);
INV_X1 g_g3904 (g3160, g3904);
INV_X1 g_g3905 (g3192, g3905);
INV_X1 g_I7517 (g3578, I7517);
INV_X1 g_g3908 (I7517, g3908);
INV_X1 g_I7520 (g2734, I7520);
INV_X1 g_g3909 (I7520, g3909);
INV_X1 g_I7523 (g2562, I7523);
INV_X1 g_g3910 (I7523, g3910);
INV_X1 g_I7526 (g2752, I7526);
INV_X1 g_g3911 (I7526, g3911);
INV_X1 g_g3912 (g3192, g3912);
INV_X1 g_g3913 (g2834, g3913);
INV_X1 g_I7545 (g3589, I7545);
INV_X1 g_g3916 (I7545, g3916);
INV_X1 g_I7548 (g3590, I7548);
INV_X1 g_g3917 (I7548, g3917);
INV_X1 g_I7551 (g2712, I7551);
INV_X1 g_g3918 (I7551, g3918);
INV_X1 g_I7554 (g2573, I7554);
INV_X1 g_g3919 (I7554, g3919);
INV_X1 g_g3920 (g3097, g3920);
INV_X1 g_I7558 (g2734, I7558);
INV_X1 g_g3921 (I7558, g3921);
INV_X1 g_I7561 (g2562, I7561);
INV_X1 g_g3922 (I7561, g3922);
INV_X1 g_I7564 (g2752, I7564);
INV_X1 g_g3923 (I7564, g3923);
INV_X1 g_I7581 (g3612, I7581);
INV_X1 g_g3926 (I7581, g3926);
INV_X1 g_I7584 (g3062, I7584);
INV_X1 g_g3927 (I7584, g3927);
INV_X1 g_g3928 (g3097, g3928);
INV_X1 g_I7588 (g2584, I7588);
INV_X1 g_g3929 (I7588, g3929);
INV_X1 g_g3930 (g3097, g3930);
INV_X1 g_I7592 (g2712, I7592);
INV_X1 g_g3931 (I7592, g3931);
INV_X1 g_I7595 (g2573, I7595);
INV_X1 g_g3932 (I7595, g3932);
INV_X1 g_g3933 (g3131, g3933);
INV_X1 g_I7599 (g2734, I7599);
INV_X1 g_g3934 (I7599, g3934);
INV_X1 g_I7602 (g2562, I7602);
INV_X1 g_g3935 (I7602, g3935);
INV_X1 g_I7605 (g2752, I7605);
INV_X1 g_g3936 (I7605, g3936);
INV_X1 g_g3937 (g2845, g3937);
INV_X1 g_I7623 (g3631, I7623);
INV_X1 g_g3940 (I7623, g3940);
INV_X1 g_I7626 (g3632, I7626);
INV_X1 g_g3941 (I7626, g3941);
INV_X1 g_I7629 (g3633, I7629);
INV_X1 g_g3942 (I7629, g3942);
INV_X1 g_I7632 (g3634, I7632);
INV_X1 g_g3943 (I7632, g3943);
INV_X1 g_I7635 (g3052, I7635);
INV_X1 g_g3944 (I7635, g3944);
INV_X1 g_g3945 (g3097, g3945);
INV_X1 g_g3946 (g3097, g3946);
INV_X1 g_I7640 (g3062, I7640);
INV_X1 g_g3947 (I7640, g3947);
INV_X1 g_g3948 (g3131, g3948);
INV_X1 g_I7644 (g2584, I7644);
INV_X1 g_g3949 (I7644, g3949);
INV_X1 g_g3950 (g3131, g3950);
INV_X1 g_I7648 (g2712, I7648);
INV_X1 g_g3951 (I7648, g3951);
INV_X1 g_I7651 (g2573, I7651);
INV_X1 g_g3952 (I7651, g3952);
INV_X1 g_g3953 (g3160, g3953);
INV_X1 g_I7655 (g2734, I7655);
INV_X1 g_g3954 (I7655, g3954);
INV_X1 g_I7658 (g2562, I7658);
INV_X1 g_g3955 (I7658, g3955);
INV_X1 g_g3956 (g2845, g3956);
INV_X1 g_I7662 (g3642, I7662);
INV_X1 g_g3957 (I7662, g3957);
INV_X1 g_g3958 (g3097, g3958);
INV_X1 g_g3959 (g3097, g3959);
INV_X1 g_I7667 (g3052, I7667);
INV_X1 g_g3960 (I7667, g3960);
INV_X1 g_g3961 (g3131, g3961);
INV_X1 g_g3962 (g3131, g3962);
INV_X1 g_I7672 (g3062, I7672);
INV_X1 g_g3963 (I7672, g3963);
INV_X1 g_g3964 (g3160, g3964);
INV_X1 g_I7676 (g2584, I7676);
INV_X1 g_g3965 (I7676, g3965);
INV_X1 g_g3966 (g3160, g3966);
INV_X1 g_I7680 (g2712, I7680);
INV_X1 g_g3967 (I7680, g3967);
INV_X1 g_I7683 (g2573, I7683);
INV_X1 g_g3968 (I7683, g3968);
INV_X1 g_g3969 (g3192, g3969);
INV_X1 g_g3970 (g2845, g3970);
INV_X1 g_I7688 (g3650, I7688);
INV_X1 g_g3971 (I7688, g3971);
INV_X1 g_I7691 (g3651, I7691);
INV_X1 g_g3972 (I7691, g3972);
INV_X1 g_g3973 (g3097, g3973);
INV_X1 g_g3974 (g3131, g3974);
INV_X1 g_g3975 (g3131, g3975);
INV_X1 g_I7697 (g3052, I7697);
INV_X1 g_g3976 (I7697, g3976);
INV_X1 g_g3977 (g3160, g3977);
INV_X1 g_g3978 (g3160, g3978);
INV_X1 g_I7702 (g3062, I7702);
INV_X1 g_g3979 (I7702, g3979);
INV_X1 g_g3980 (g3192, g3980);
INV_X1 g_I7706 (g2584, I7706);
INV_X1 g_g3981 (I7706, g3981);
INV_X1 g_g3982 (g3192, g3982);
INV_X1 g_g3983 (g2845, g3983);
INV_X1 g_I7712 (g3657, I7712);
INV_X1 g_g3985 (I7712, g3985);
INV_X1 g_I7716 (g3038, I7716);
INV_X1 g_g3987 (I7716, g3987);
INV_X1 g_g3988 (g3097, g3988);
INV_X1 g_g3989 (g3131, g3989);
INV_X1 g_g3990 (g3160, g3990);
INV_X1 g_g3991 (g3160, g3991);
INV_X1 g_I7723 (g3052, I7723);
INV_X1 g_g3992 (I7723, g3992);
INV_X1 g_g3993 (g3192, g3993);
INV_X1 g_g3994 (g3192, g3994);
INV_X1 g_I7728 (g3675, I7728);
INV_X1 g_g3995 (I7728, g3995);
INV_X1 g_I7731 (g3029, I7731);
INV_X1 g_g3996 (I7731, g3996);
INV_X1 g_I7734 (g2595, I7734);
INV_X1 g_g3997 (I7734, g3997);
INV_X1 g_g3998 (g3097, g3998);
INV_X1 g_I7738 (g3038, I7738);
INV_X1 g_g3999 (I7738, g3999);
INV_X1 g_g4000 (g3131, g4000);
INV_X1 g_g4001 (g3160, g4001);
INV_X1 g_g4002 (g3192, g4002);
INV_X1 g_g4003 (g3192, g4003);
INV_X1 g_g4004 (g2845, g4004);
INV_X1 g_I7746 (g3591, I7746);
INV_X1 g_g4005 (I7746, g4005);
INV_X1 g_I7749 (g3692, I7749);
INV_X1 g_g4006 (I7749, g4006);
INV_X1 g_I7752 (g3591, I7752);
INV_X1 g_g4007 (I7752, g4007);
INV_X1 g_I7755 (g3019, I7755);
INV_X1 g_g4008 (I7755, g4008);
INV_X1 g_I7758 (g2605, I7758);
INV_X1 g_g4009 (I7758, g4009);
INV_X1 g_g4010 (g3097, g4010);
INV_X1 g_I7762 (g3029, I7762);
INV_X1 g_g4011 (I7762, g4011);
INV_X1 g_I7765 (g2595, I7765);
INV_X1 g_g4012 (I7765, g4012);
INV_X1 g_g4013 (g3131, g4013);
INV_X1 g_I7769 (g3038, I7769);
INV_X1 g_g4014 (I7769, g4014);
INV_X1 g_g4015 (g3160, g4015);
INV_X1 g_g4016 (g3192, g4016);
INV_X1 g_g4017 (g2845, g4017);
INV_X1 g_I7775 (g3705, I7775);
INV_X1 g_g4018 (I7775, g4018);
INV_X1 g_I7778 (g3019, I7778);
INV_X1 g_g4019 (I7778, g4019);
INV_X1 g_I7781 (g2605, I7781);
INV_X1 g_g4020 (I7781, g4020);
INV_X1 g_g4021 (g3131, g4021);
INV_X1 g_I7785 (g3029, I7785);
INV_X1 g_g4022 (I7785, g4022);
INV_X1 g_I7788 (g2595, I7788);
INV_X1 g_g4023 (I7788, g4023);
INV_X1 g_g4024 (g3160, g4024);
INV_X1 g_I7792 (g3038, I7792);
INV_X1 g_g4025 (I7792, g4025);
INV_X1 g_g4026 (g3192, g4026);
INV_X1 g_g4027 (g2845, g4027);
INV_X1 g_I7797 (g3019, I7797);
INV_X1 g_g4028 (I7797, g4028);
INV_X1 g_I7800 (g2605, I7800);
INV_X1 g_g4029 (I7800, g4029);
INV_X1 g_g4030 (g3160, g4030);
INV_X1 g_I7804 (g3029, I7804);
INV_X1 g_g4031 (I7804, g4031);
INV_X1 g_I7807 (g2595, I7807);
INV_X1 g_g4032 (I7807, g4032);
INV_X1 g_g4033 (g3192, g4033);
INV_X1 g_I7811 (g3019, I7811);
INV_X1 g_g4034 (I7811, g4034);
INV_X1 g_I7814 (g2605, I7814);
INV_X1 g_g4035 (I7814, g4035);
INV_X1 g_g4036 (g3192, g4036);
INV_X1 g_g4037 (g2845, g4037);
INV_X1 g_g4041 (g2605, g4041);
INV_X1 g_g4044 (g2595, g4044);
INV_X1 g_g4050 (g3080, g4050);
INV_X1 g_g4051 (g3093, g4051);
INV_X1 g_g4056 (g3082, g4056);
INV_X1 g_I7832 (g2768, I7832);
INV_X1 g_g4057 (I7832, g4057);
INV_X1 g_I7838 (g2781, I7838);
INV_X1 g_g4065 (I7838, g4065);
INV_X1 g_I7844 (g3784, I7844);
INV_X1 g_g4069 (I7844, g4069);
INV_X1 g_I7847 (g3798, I7847);
INV_X1 g_g4070 (I7847, g4070);
INV_X1 g_I7850 (g2795, I7850);
INV_X1 g_g4071 (I7850, g4071);
INV_X1 g_I7856 (g3805, I7856);
INV_X1 g_g4075 (I7856, g4075);
INV_X1 g_I7859 (g2804, I7859);
INV_X1 g_g4076 (I7859, g4076);
INV_X1 g_I7864 (g3812, I7864);
INV_X1 g_g4079 (I7864, g4079);
INV_X1 g_I7867 (g2818, I7867);
INV_X1 g_g4080 (I7867, g4080);
INV_X1 g_I7870 (g2827, I7870);
INV_X1 g_g4081 (I7870, g4081);
INV_X1 g_I7875 (g3819, I7875);
INV_X1 g_g4084 (I7875, g4084);
INV_X1 g_I7878 (g2829, I7878);
INV_X1 g_g4085 (I7878, g4085);
INV_X1 g_I7882 (g2700, I7882);
INV_X1 g_g4087 (I7882, g4087);
INV_X1 g_I7885 (g2837, I7885);
INV_X1 g_g4088 (I7885, g4088);
INV_X1 g_I7888 (g3505, I7888);
INV_X1 g_g4089 (I7888, g4089);
INV_X1 g_I7899 (g3743, I7899);
INV_X1 g_g4092 (I7899, g4092);
INV_X1 g_I7902 (g2709, I7902);
INV_X1 g_g4093 (I7902, g4093);
INV_X1 g_I7905 (g2863, I7905);
INV_X1 g_g4094 (I7905, g4094);
INV_X1 g_I7908 (g3516, I7908);
INV_X1 g_g4095 (I7908, g4095);
INV_X1 g_I7911 (g2767, I7911);
INV_X1 g_g4096 (I7911, g4096);
INV_X1 g_I7919 (g3761, I7919);
INV_X1 g_g4102 (I7919, g4102);
INV_X1 g_I7922 (g3462, I7922);
INV_X1 g_g4103 (I7922, g4103);
INV_X1 g_I7925 (g2761, I7925);
INV_X1 g_g4104 (I7925, g4104);
INV_X1 g_I7928 (g2873, I7928);
INV_X1 g_g4105 (I7928, g4105);
INV_X1 g_I7931 (g2780, I7931);
INV_X1 g_g4106 (I7931, g4106);
INV_X1 g_I7944 (g3774, I7944);
INV_X1 g_g4111 (I7944, g4111);
INV_X1 g_I7947 (g3485, I7947);
INV_X1 g_g4112 (I7947, g4112);
INV_X1 g_I7950 (g2774, I7950);
INV_X1 g_g4113 (I7950, g4113);
INV_X1 g_I7953 (g3542, I7953);
INV_X1 g_g4114 (I7953, g4114);
INV_X1 g_I7956 (g2810, I7956);
INV_X1 g_g4115 (I7956, g4115);
INV_X1 g_I7959 (g2793, I7959);
INV_X1 g_g4116 (I7959, g4116);
INV_X1 g_I7964 (g3488, I7964);
INV_X1 g_g4119 (I7964, g4119);
INV_X1 g_I7967 (g2787, I7967);
INV_X1 g_g4120 (I7967, g4120);
INV_X1 g_I7970 (g3557, I7970);
INV_X1 g_g4121 (I7970, g4121);
INV_X1 g_I7973 (g3071, I7973);
INV_X1 g_g4122 (I7973, g4122);
INV_X1 g_I7978 (g3574, I7978);
INV_X1 g_g4125 (I7978, g4125);
INV_X1 g_I7981 (g3555, I7981);
INV_X1 g_g4126 (I7981, g4126);
INV_X1 g_I7987 (g3528, I7987);
INV_X1 g_g4130 (I7987, g4130);
INV_X1 g_g4134 (g3676, g4134);
INV_X1 g_I8011 (g3225, I8011);
INV_X1 g_g4146 (I8011, g4146);
INV_X1 g_I8024 (g3076, I8024);
INV_X1 g_g4153 (I8024, g4153);
INV_X1 g_I8084 (g3706, I8084);
INV_X1 g_g4191 (I8084, g4191);
INV_X1 g_I8094 (g2976, I8094);
INV_X1 g_g4195 (I8094, g4195);
INV_X1 g_I8097 (g3237, I8097);
INV_X1 g_g4196 (I8097, g4196);
INV_X1 g_g4197 (g3591, g4197);
INV_X1 g_I8101 (g3259, I8101);
INV_X1 g_g4198 (I8101, g4198);
INV_X1 g_I8105 (g3339, I8105);
INV_X1 g_g4200 (I8105, g4200);
INV_X1 g_g4202 (g2810, g4202);
INV_X1 g_g4226 (g3591, g4226);
INV_X1 g_I8140 (g3429, I8140);
INV_X1 g_g4229 (I8140, g4229);
INV_X1 g_I8161 (g3517, I8161);
INV_X1 g_g4242 (I8161, g4242);
INV_X1 g_I8172 (g3524, I8172);
INV_X1 g_g4245 (I8172, g4245);
INV_X1 g_I8177 (g2810, I8177);
INV_X1 g_g4250 (I8177, g4250);
INV_X1 g_I8180 (g3529, I8180);
INV_X1 g_g4251 (I8180, g4251);
INV_X1 g_g4253 (g2734, g4253);
INV_X1 g_I8190 (g3545, I8190);
INV_X1 g_g4257 (I8190, g4257);
INV_X1 g_I8193 (g3547, I8193);
INV_X1 g_g4258 (I8193, g4258);
INV_X1 g_I8196 (g3654, I8196);
INV_X1 g_g4259 (I8196, g4259);
INV_X1 g_g4265 (g3591, g4265);
INV_X1 g_I8202 (g3560, I8202);
INV_X1 g_g4266 (I8202, g4266);
INV_X1 g_I8205 (g2655, I8205);
INV_X1 g_g4267 (I8205, g4267);
INV_X1 g_g4270 (g2573, g4270);
INV_X1 g_I8215 (g3577, I8215);
INV_X1 g_g4273 (I8215, g4273);
INV_X1 g_I8218 (g3002, I8218);
INV_X1 g_g4274 (I8218, g4274);
INV_X1 g_g4275 (g3790, g4275);
INV_X1 g_g4279 (g3340, g4279);
INV_X1 g_g4281 (g2562, g4281);
INV_X1 g_I8233 (g3588, I8233);
INV_X1 g_g4285 (I8233, g4285);
INV_X1 g_g4286 (g3790, g4286);
INV_X1 g_g4296 (g3790, g4296);
INV_X1 g_I8261 (g3643, I8261);
INV_X1 g_g4300 (I8261, g4300);
INV_X1 g_I8264 (g3653, I8264);
INV_X1 g_g4301 (I8264, g4301);
INV_X1 g_I8268 (g2801, I8268);
INV_X1 g_g4303 (I8268, g4303);
INV_X1 g_I8273 (g2976, I8273);
INV_X1 g_g4306 (I8273, g4306);
INV_X1 g_g4307 (g3700, g4307);
INV_X1 g_I8277 (g3504, I8277);
INV_X1 g_g4308 (I8277, g4308);
INV_X1 g_I8282 (g3515, I8282);
INV_X1 g_g4311 (I8282, g4311);
INV_X1 g_I8291 (g878, I8291);
INV_X1 g_g4316 (I8291, g4316);
INV_X1 g_g4328 (g3086, g4328);
INV_X1 g_g4335 (g3659, g4335);
INV_X1 g_I8308 (g3674, I8308);
INV_X1 g_g4341 (I8308, g4341);
INV_X1 g_g4344 (g3124, g4344);
INV_X1 g_I8315 (g3691, I8315);
INV_X1 g_g4350 (I8315, g4350);
INV_X1 g_g4353 (g3665, g4353);
INV_X1 g_g4357 (g3679, g4357);
INV_X1 g_g4358 (g3680, g4358);
INV_X1 g_I8333 (g3721, I8333);
INV_X1 g_g4360 (I8333, g4360);
INV_X1 g_g4362 (g2810, g4362);
INV_X1 g_I8351 (g1160, I8351);
INV_X1 g_g4370 (I8351, g4370);
INV_X1 g_I8354 (g1163, I8354);
INV_X1 g_g4371 (I8354, g4371);
INV_X1 g_I8357 (g1182, I8357);
INV_X1 g_g4372 (I8357, g4372);
INV_X1 g_I8360 (g1186, I8360);
INV_X1 g_g4373 (I8360, g4373);
INV_X1 g_g4381 (g3466, g4381);
INV_X1 g_I8373 (g3783, I8373);
INV_X1 g_g4382 (I8373, g4382);
INV_X1 g_I8428 (g3611, I8428);
INV_X1 g_g4426 (I8428, g4426);
INV_X1 g_I8446 (g3014, I8446);
INV_X1 g_g4438 (I8446, g4438);
INV_X1 g_I8449 (g3630, I8449);
INV_X1 g_g4443 (I8449, g4443);
INV_X1 g_I8452 (g2816, I8452);
INV_X1 g_g4444 (I8452, g4444);
INV_X1 g_g4455 (g3811, g4455);
INV_X1 g_I8477 (g3014, I8477);
INV_X1 g_g4457 (I8477, g4457);
INV_X1 g_I8480 (g3640, I8480);
INV_X1 g_g4462 (I8480, g4462);
INV_X1 g_I8483 (g3641, I8483);
INV_X1 g_g4463 (I8483, g4463);
INV_X1 g_I8486 (g2824, I8486);
INV_X1 g_g4464 (I8486, g4464);
INV_X1 g_g4465 (g3677, g4465);
INV_X1 g_g4475 (g3818, g4475);
INV_X1 g_I8517 (g3014, I8517);
INV_X1 g_g4477 (I8517, g4477);
INV_X1 g_I8520 (g3652, I8520);
INV_X1 g_g4482 (I8520, g4482);
INV_X1 g_g4489 (g2826, g4489);
INV_X1 g_I8543 (g2810, I8543);
INV_X1 g_g4493 (I8543, g4493);
INV_X1 g_g4500 (g2832, g4500);
INV_X1 g_g4501 (g2801, g4501);
INV_X1 g_I8565 (g3071, I8565);
INV_X1 g_g4503 (I8565, g4503);
INV_X1 g_g4510 (g2840, g4510);
INV_X1 g_g4511 (g2841, g4511);
INV_X1 g_g4512 (g2842, g4512);
INV_X1 g_g4521 (g2866, g4521);
INV_X1 g_g4522 (g2867, g4522);
INV_X1 g_g4523 (g2868, g4523);
INV_X1 g_g4524 (g2869, g4524);
INV_X1 g_g4525 (g2870, g4525);
INV_X1 g_g4527 (g3466, g4527);
INV_X1 g_g4535 (g2876, g4535);
INV_X1 g_g4536 (g2877, g4536);
INV_X1 g_g4537 (g2878, g4537);
INV_X1 g_g4538 (g2880, g4538);
INV_X1 g_g4539 (g2881, g4539);
INV_X1 g_g4540 (g2882, g4540);
INV_X1 g_g4541 (g2883, g4541);
INV_X1 g_g4542 (g2884, g4542);
INV_X1 g_g4543 (g2885, g4543);
INV_X1 g_g4544 (g2886, g4544);
INV_X1 g_g4545 (g2887, g4545);
INV_X1 g_g4547 (g3466, g4547);
INV_X1 g_g4552 (g2890, g4552);
INV_X1 g_g4553 (g2891, g4553);
INV_X1 g_g4554 (g2892, g4554);
INV_X1 g_g4555 (g2894, g4555);
INV_X1 g_g4556 (g2895, g4556);
INV_X1 g_g4557 (g2896, g4557);
INV_X1 g_g4558 (g2897, g4558);
INV_X1 g_g4559 (g2898, g4559);
INV_X1 g_g4560 (g2899, g4560);
INV_X1 g_g4561 (g2900, g4561);
INV_X1 g_g4562 (g3466, g4562);
INV_X1 g_I8665 (g3051, I8665);
INV_X1 g_g4564 (I8665, g4564);
INV_X1 g_g4565 (g2901, g4565);
INV_X1 g_g4566 (g2902, g4566);
INV_X1 g_g4567 (g2903, g4567);
INV_X1 g_g4568 (g2904, g4568);
INV_X1 g_g4569 (g2906, g4569);
INV_X1 g_g4570 (g2907, g4570);
INV_X1 g_g4571 (g2908, g4571);
INV_X1 g_g4572 (g2909, g4572);
INV_X1 g_g4573 (g2911, g4573);
INV_X1 g_g4574 (g3466, g4574);
INV_X1 g_g4576 (g2913, g4576);
INV_X1 g_g4577 (g2914, g4577);
INV_X1 g_g4578 (g2917, g4578);
INV_X1 g_g4579 (g2918, g4579);
INV_X1 g_g4580 (g2919, g4580);
INV_X1 g_g4581 (g2921, g4581);
INV_X1 g_g4582 (g2922, g4582);
INV_X1 g_g4583 (g2924, g4583);
INV_X1 g_g4584 (g3466, g4584);
INV_X1 g_g4585 (g2925, g4585);
INV_X1 g_g4586 (g2926, g4586);
INV_X1 g_g4587 (g2928, g4587);
INV_X1 g_g4588 (g2929, g4588);
INV_X1 g_g4589 (g2930, g4589);
INV_X1 g_g4590 (g2932, g4590);
INV_X1 g_g4591 (g2937, g4591);
INV_X1 g_g4592 (g2938, g4592);
INV_X1 g_g4593 (g2939, g4593);
INV_X1 g_g4594 (g2941, g4594);
INV_X1 g_g4595 (g2942, g4595);
INV_X1 g_g4596 (g3466, g4596);
INV_X1 g_I8706 (g3828, I8706);
INV_X1 g_g4597 (I8706, g4597);
INV_X1 g_I8709 (g4191, I8709);
INV_X1 g_g4598 (I8709, g4598);
INV_X1 g_I8712 (g4007, I8712);
INV_X1 g_g4599 (I8712, g4599);
INV_X1 g_I8715 (g3903, I8715);
INV_X1 g_g4600 (I8715, g4600);
INV_X1 g_I8718 (g3909, I8718);
INV_X1 g_g4601 (I8718, g4601);
INV_X1 g_I8721 (g3918, I8721);
INV_X1 g_g4602 (I8721, g4602);
INV_X1 g_I8724 (g3927, I8724);
INV_X1 g_g4603 (I8724, g4603);
INV_X1 g_I8727 (g3944, I8727);
INV_X1 g_g4604 (I8727, g4604);
INV_X1 g_I8730 (g3987, I8730);
INV_X1 g_g4605 (I8730, g4605);
INV_X1 g_I8733 (g3996, I8733);
INV_X1 g_g4606 (I8733, g4606);
INV_X1 g_I8736 (g4008, I8736);
INV_X1 g_g4607 (I8736, g4607);
INV_X1 g_I8739 (g3910, I8739);
INV_X1 g_g4608 (I8739, g4608);
INV_X1 g_I8742 (g3919, I8742);
INV_X1 g_g4609 (I8742, g4609);
INV_X1 g_I8745 (g3929, I8745);
INV_X1 g_g4610 (I8745, g4610);
INV_X1 g_I8748 (g3997, I8748);
INV_X1 g_g4611 (I8748, g4611);
INV_X1 g_I8751 (g4009, I8751);
INV_X1 g_g4612 (I8751, g4612);
INV_X1 g_I8754 (g3911, I8754);
INV_X1 g_g4613 (I8754, g4613);
INV_X1 g_I8757 (g3921, I8757);
INV_X1 g_g4614 (I8757, g4614);
INV_X1 g_I8760 (g3931, I8760);
INV_X1 g_g4615 (I8760, g4615);
INV_X1 g_I8763 (g3947, I8763);
INV_X1 g_g4616 (I8763, g4616);
INV_X1 g_I8766 (g3960, I8766);
INV_X1 g_g4617 (I8766, g4617);
INV_X1 g_I8769 (g3999, I8769);
INV_X1 g_g4618 (I8769, g4618);
INV_X1 g_I8772 (g4011, I8772);
INV_X1 g_g4619 (I8772, g4619);
INV_X1 g_I8775 (g4019, I8775);
INV_X1 g_g4620 (I8775, g4620);
INV_X1 g_I8778 (g3922, I8778);
INV_X1 g_g4621 (I8778, g4621);
INV_X1 g_I8781 (g3932, I8781);
INV_X1 g_g4622 (I8781, g4622);
INV_X1 g_I8784 (g3949, I8784);
INV_X1 g_g4623 (I8784, g4623);
INV_X1 g_I8787 (g4012, I8787);
INV_X1 g_g4624 (I8787, g4624);
INV_X1 g_I8790 (g4020, I8790);
INV_X1 g_g4625 (I8790, g4625);
INV_X1 g_I8793 (g3923, I8793);
INV_X1 g_g4626 (I8793, g4626);
INV_X1 g_I8796 (g3934, I8796);
INV_X1 g_g4627 (I8796, g4627);
INV_X1 g_I8799 (g3951, I8799);
INV_X1 g_g4628 (I8799, g4628);
INV_X1 g_I8802 (g3963, I8802);
INV_X1 g_g4629 (I8802, g4629);
INV_X1 g_I8805 (g3976, I8805);
INV_X1 g_g4630 (I8805, g4630);
INV_X1 g_I8808 (g4014, I8808);
INV_X1 g_g4631 (I8808, g4631);
INV_X1 g_I8811 (g4022, I8811);
INV_X1 g_g4632 (I8811, g4632);
INV_X1 g_I8814 (g4028, I8814);
INV_X1 g_g4633 (I8814, g4633);
INV_X1 g_I8817 (g3935, I8817);
INV_X1 g_g4634 (I8817, g4634);
INV_X1 g_I8820 (g3952, I8820);
INV_X1 g_g4635 (I8820, g4635);
INV_X1 g_I8823 (g3965, I8823);
INV_X1 g_g4636 (I8823, g4636);
INV_X1 g_I8826 (g4023, I8826);
INV_X1 g_g4637 (I8826, g4637);
INV_X1 g_I8829 (g4029, I8829);
INV_X1 g_g4638 (I8829, g4638);
INV_X1 g_I8832 (g3936, I8832);
INV_X1 g_g4639 (I8832, g4639);
INV_X1 g_I8835 (g3954, I8835);
INV_X1 g_g4640 (I8835, g4640);
INV_X1 g_I8838 (g3967, I8838);
INV_X1 g_g4641 (I8838, g4641);
INV_X1 g_I8841 (g3979, I8841);
INV_X1 g_g4642 (I8841, g4642);
INV_X1 g_I8844 (g3992, I8844);
INV_X1 g_g4643 (I8844, g4643);
INV_X1 g_I8847 (g4025, I8847);
INV_X1 g_g4644 (I8847, g4644);
INV_X1 g_I8850 (g4031, I8850);
INV_X1 g_g4645 (I8850, g4645);
INV_X1 g_I8853 (g4034, I8853);
INV_X1 g_g4646 (I8853, g4646);
INV_X1 g_I8856 (g3955, I8856);
INV_X1 g_g4647 (I8856, g4647);
INV_X1 g_I8859 (g3968, I8859);
INV_X1 g_g4648 (I8859, g4648);
INV_X1 g_I8862 (g3981, I8862);
INV_X1 g_g4649 (I8862, g4649);
INV_X1 g_I8865 (g4032, I8865);
INV_X1 g_g4650 (I8865, g4650);
INV_X1 g_I8868 (g4035, I8868);
INV_X1 g_g4651 (I8868, g4651);
INV_X1 g_I8871 (g3869, I8871);
INV_X1 g_g4652 (I8871, g4652);
INV_X1 g_I8874 (g3884, I8874);
INV_X1 g_g4653 (I8874, g4653);
INV_X1 g_I8877 (g4274, I8877);
INV_X1 g_g4654 (I8877, g4654);
INV_X1 g_I8880 (g4303, I8880);
INV_X1 g_g4655 (I8880, g4655);
INV_X1 g_I8883 (g4198, I8883);
INV_X1 g_g4656 (I8883, g4656);
INV_X1 g_I8886 (g4308, I8886);
INV_X1 g_g4657 (I8886, g4657);
INV_X1 g_I8889 (g4311, I8889);
INV_X1 g_g4658 (I8889, g4658);
INV_X1 g_I8892 (g4115, I8892);
INV_X1 g_g4659 (I8892, g4659);
INV_X1 g_I8895 (g4130, I8895);
INV_X1 g_g4660 (I8895, g4660);
INV_X1 g_I8898 (g4089, I8898);
INV_X1 g_g4661 (I8898, g4661);
INV_X1 g_I8901 (g4122, I8901);
INV_X1 g_g4662 (I8901, g4662);
INV_X1 g_I8904 (g4126, I8904);
INV_X1 g_g4663 (I8904, g4663);
INV_X1 g_I8907 (g4095, I8907);
INV_X1 g_g4664 (I8907, g4664);
INV_X1 g_I8910 (g4200, I8910);
INV_X1 g_g4665 (I8910, g4665);
INV_X1 g_I8913 (g4306, I8913);
INV_X1 g_g4666 (I8913, g4666);
INV_X1 g_I8916 (g4195, I8916);
INV_X1 g_g4667 (I8916, g4667);
INV_X1 g_I8919 (g4196, I8919);
INV_X1 g_g4668 (I8919, g4668);
INV_X1 g_I8922 (g4229, I8922);
INV_X1 g_g4669 (I8922, g4669);
INV_X1 g_I8925 (g4482, I8925);
INV_X1 g_g4670 (I8925, g4670);
INV_X1 g_I8928 (g4153, I8928);
INV_X1 g_g4673 (I8928, g4673);
INV_X1 g_I8932 (g4096, I8932);
INV_X1 g_g4677 (I8932, g4677);
INV_X1 g_I8935 (g4005, I8935);
INV_X1 g_g4678 (I8935, g4678);
INV_X1 g_I8945 (g4106, I8945);
INV_X1 g_g4680 (I8945, g4680);
INV_X1 g_I8949 (g4116, I8949);
INV_X1 g_g4684 (I8949, g4684);
INV_X1 g_I8952 (g4197, I8952);
INV_X1 g_g4685 (I8952, g4685);
INV_X1 g_I8962 (g4553, I8962);
INV_X1 g_g4687 (I8962, g4687);
INV_X1 g_I8966 (g4444, I8966);
INV_X1 g_g4689 (I8966, g4689);
INV_X1 g_I8971 (g4464, I8971);
INV_X1 g_g4692 (I8971, g4692);
INV_X1 g_I8974 (g3871, I8974);
INV_X1 g_g4693 (I8974, g4693);
INV_X1 g_I8977 (g3877, I8977);
INV_X1 g_g4694 (I8977, g4694);
INV_X1 g_I8980 (g4535, I8980);
INV_X1 g_g4695 (I8980, g4695);
INV_X1 g_I8983 (g4536, I8983);
INV_X1 g_g4696 (I8983, g4696);
INV_X1 g_I8986 (g4552, I8986);
INV_X1 g_g4697 (I8986, g4697);
INV_X1 g_I8989 (g4537, I8989);
INV_X1 g_g4698 (I8989, g4698);
INV_X1 g_I8994 (g4565, I8994);
INV_X1 g_g4701 (I8994, g4701);
INV_X1 g_I8998 (g4576, I8998);
INV_X1 g_g4703 (I8998, g4703);
INV_X1 g_I9001 (g4577, I9001);
INV_X1 g_g4704 (I9001, g4704);
INV_X1 g_I9005 (g4585, I9005);
INV_X1 g_g4706 (I9005, g4706);
INV_X1 g_I9009 (g4591, I9009);
INV_X1 g_g4710 (I9009, g4710);
INV_X1 g_I9014 (g3864, I9014);
INV_X1 g_g4713 (I9014, g4713);
INV_X1 g_I9018 (g3872, I9018);
INV_X1 g_g4718 (I9018, g4718);
INV_X1 g_I9021 (g4489, I9021);
INV_X1 g_g4719 (I9021, g4719);
INV_X1 g_I9025 (g4462, I9025);
INV_X1 g_g4721 (I9025, g4721);
INV_X1 g_I9034 (g4317, I9034);
INV_X1 g_g4732 (I9034, g4732);
INV_X1 g_g4733 (g4202, g4733);
INV_X1 g_I9050 (g3881, I9050);
INV_X1 g_g4738 (I9050, g4738);
INV_X1 g_I9053 (g4327, I9053);
INV_X1 g_g4739 (I9053, g4739);
INV_X1 g_I9064 (g4302, I9064);
INV_X1 g_g4742 (I9064, g4742);
INV_X1 g_I9076 (g4353, I9076);
INV_X1 g_g4746 (I9076, g4746);
INV_X1 g_g4748 (g4465, g4748);
INV_X1 g_I9081 (g4357, I9081);
INV_X1 g_g4776 (I9081, g4776);
INV_X1 g_I9084 (g4358, I9084);
INV_X1 g_g4777 (I9084, g4777);
INV_X1 g_I9089 (g4566, I9089);
INV_X1 g_g4780 (I9089, g4780);
INV_X1 g_I9095 (g4283, I9095);
INV_X1 g_g4784 (I9095, g4784);
INV_X1 g_I9103 (g4374, I9103);
INV_X1 g_g4788 (I9103, g4788);
INV_X1 g_I9111 (g4232, I9111);
INV_X1 g_g4792 (I9111, g4792);
INV_X1 g_I9116 (g4297, I9116);
INV_X1 g_g4795 (I9116, g4795);
INV_X1 g_I9123 (g4455, I9123);
INV_X1 g_g4800 (I9123, g4800);
INV_X1 g_I9126 (g3870, I9126);
INV_X1 g_g4801 (I9126, g4801);
INV_X1 g_I9129 (g4475, I9129);
INV_X1 g_g4802 (I9129, g4802);
INV_X1 g_I9132 (g4284, I9132);
INV_X1 g_g4803 (I9132, g4803);
INV_X1 g_I9136 (g4280, I9136);
INV_X1 g_g4805 (I9136, g4805);
INV_X1 g_I9139 (g4364, I9139);
INV_X1 g_g4806 (I9139, g4806);
INV_X1 g_I9142 (g4236, I9142);
INV_X1 g_g4807 (I9142, g4807);
INV_X1 g_I9145 (g4264, I9145);
INV_X1 g_g4808 (I9145, g4808);
INV_X1 g_I9148 (g4354, I9148);
INV_X1 g_g4809 (I9148, g4809);
INV_X1 g_I9158 (g4256, I9158);
INV_X1 g_g4811 (I9158, g4811);
INV_X1 g_I9162 (g4272, I9162);
INV_X1 g_g4813 (I9162, g4813);
INV_X1 g_I9177 (g4299, I9177);
INV_X1 g_g4822 (I9177, g4822);
INV_X1 g_g4841 (g4250, g4841);
INV_X1 g_I9209 (g4349, I9209);
INV_X1 g_g4867 (I9209, g4867);
INV_X1 g_I9217 (g4443, I9217);
INV_X1 g_g4873 (I9217, g4873);
INV_X1 g_g4882 (g4069, g4882);
INV_X1 g_g4885 (g4070, g4885);
INV_X1 g_g4886 (g4071, g4886);
INV_X1 g_g4890 (g4075, g4890);
INV_X1 g_g4891 (g4076, g4891);
INV_X1 g_I9250 (g4134, I9250);
INV_X1 g_g4892 (I9250, g4892);
INV_X1 g_g4895 (g4078, g4895);
INV_X1 g_g4898 (g4079, g4898);
INV_X1 g_g4899 (g4080, g4899);
INV_X1 g_I9258 (g4249, I9258);
INV_X1 g_g4900 (I9258, g4900);
INV_X1 g_g4903 (g4084, g4903);
INV_X1 g_g4904 (g4085, g4904);
INV_X1 g_g4907 (g4087, g4907);
INV_X1 g_g4908 (g4088, g4908);
INV_X1 g_I9271 (g4263, I9271);
INV_X1 g_g4909 (I9271, g4909);
INV_X1 g_g4913 (g4092, g4913);
INV_X1 g_g4914 (g4093, g4914);
INV_X1 g_g4915 (g4094, g4915);
INV_X1 g_g4916 (g4202, g4916);
INV_X1 g_g4917 (g4102, g4917);
INV_X1 g_g4918 (g4103, g4918);
INV_X1 g_g4919 (g4104, g4919);
INV_X1 g_g4920 (g4105, g4920);
INV_X1 g_g4921 (g4202, g4921);
INV_X1 g_g4922 (g4111, g4922);
INV_X1 g_g4923 (g4112, g4923);
INV_X1 g_g4924 (g4113, g4924);
INV_X1 g_g4925 (g4114, g4925);
INV_X1 g_g4926 (g4202, g4926);
INV_X1 g_g4928 (g4119, g4928);
INV_X1 g_g4929 (g4120, g4929);
INV_X1 g_g4930 (g4121, g4930);
INV_X1 g_I9301 (g4295, I9301);
INV_X1 g_g4931 (I9301, g4931);
INV_X1 g_g4932 (g4202, g4932);
INV_X1 g_g4934 (g4125, g4934);
INV_X1 g_g4935 (g4202, g4935);
INV_X1 g_I9310 (g4268, I9310);
INV_X1 g_g4938 (I9310, g4938);
INV_X1 g_g4960 (g4259, g4960);
INV_X1 g_g4963 (g4328, g4963);
INV_X1 g_I9325 (g4242, I9325);
INV_X1 g_g5000 (I9325, g5000);
INV_X1 g_g5002 (g4335, g5002);
INV_X1 g_I9333 (g4245, I9333);
INV_X1 g_g5006 (I9333, g5006);
INV_X1 g_I9336 (g4493, I9336);
INV_X1 g_g5007 (I9336, g5007);
INV_X1 g_g5009 (g4344, g5009);
INV_X1 g_I9341 (g4251, I9341);
INV_X1 g_g5013 (I9341, g5013);
INV_X1 g_I9344 (g4341, I9344);
INV_X1 g_g5014 (I9344, g5014);
INV_X1 g_I9347 (g3896, I9347);
INV_X1 g_g5015 (I9347, g5015);
INV_X1 g_I9350 (g4503, I9350);
INV_X1 g_g5016 (I9350, g5016);
INV_X1 g_g5022 (g4438, g5022);
INV_X1 g_I9360 (g4257, I9360);
INV_X1 g_g5024 (I9360, g5024);
INV_X1 g_I9363 (g4258, I9363);
INV_X1 g_g5025 (I9363, g5025);
INV_X1 g_I9366 (g4350, I9366);
INV_X1 g_g5026 (I9366, g5026);
INV_X1 g_I9369 (g3901, I9369);
INV_X1 g_g5027 (I9369, g5027);
INV_X1 g_I9372 (g3902, I9372);
INV_X1 g_g5028 (I9372, g5028);
INV_X1 g_g5037 (g4438, g5037);
INV_X1 g_g5038 (g4457, g5038);
INV_X1 g_I9393 (g4266, I9393);
INV_X1 g_g5041 (I9393, g5041);
INV_X1 g_I9396 (g3908, I9396);
INV_X1 g_g5042 (I9396, g5042);
INV_X1 g_I9407 (g4232, I9407);
INV_X1 g_g5051 (I9407, g5051);
INV_X1 g_g5053 (g4438, g5053);
INV_X1 g_g5054 (g4457, g5054);
INV_X1 g_g5055 (g4477, g5055);
INV_X1 g_I9416 (g4273, I9416);
INV_X1 g_g5058 (I9416, g5058);
INV_X1 g_I9419 (g3916, I9419);
INV_X1 g_g5059 (I9419, g5059);
INV_X1 g_I9422 (g4360, I9422);
INV_X1 g_g5060 (I9422, g5060);
INV_X1 g_I9425 (g3917, I9425);
INV_X1 g_g5061 (I9425, g5061);
INV_X1 g_g5071 (g4438, g5071);
INV_X1 g_g5072 (g4457, g5072);
INV_X1 g_g5073 (g4477, g5073);
INV_X1 g_I9440 (g4285, I9440);
INV_X1 g_g5074 (I9440, g5074);
INV_X1 g_I9443 (g4564, I9443);
INV_X1 g_g5075 (I9443, g5075);
INV_X1 g_I9446 (g3926, I9446);
INV_X1 g_g5076 (I9446, g5076);
INV_X1 g_g5083 (g4457, g5083);
INV_X1 g_g5084 (g4477, g5084);
INV_X1 g_I9457 (g3940, I9457);
INV_X1 g_g5085 (I9457, g5085);
INV_X1 g_I9460 (g3941, I9460);
INV_X1 g_g5086 (I9460, g5086);
INV_X1 g_I9463 (g3942, I9463);
INV_X1 g_g5087 (I9463, g5087);
INV_X1 g_I9466 (g3943, I9466);
INV_X1 g_g5088 (I9466, g5088);
INV_X1 g_g5099 (g4477, g5099);
INV_X1 g_I9484 (g3957, I9484);
INV_X1 g_g5100 (I9484, g5100);
INV_X1 g_g5101 (g4259, g5101);
INV_X1 g_I9493 (g4426, I9493);
INV_X1 g_g5109 (I9493, g5109);
INV_X1 g_I9496 (g3971, I9496);
INV_X1 g_g5112 (I9496, g5112);
INV_X1 g_I9499 (g4382, I9499);
INV_X1 g_g5113 (I9499, g5113);
INV_X1 g_I9502 (g3972, I9502);
INV_X1 g_g5114 (I9502, g5114);
INV_X1 g_I9505 (g4300, I9505);
INV_X1 g_g5115 (I9505, g5115);
INV_X1 g_I9512 (g3985, I9512);
INV_X1 g_g5120 (I9512, g5120);
INV_X1 g_I9515 (g4301, I9515);
INV_X1 g_g5121 (I9515, g5121);
INV_X1 g_I9520 (g3995, I9520);
INV_X1 g_g5124 (I9520, g5124);
INV_X1 g_I9525 (g4413, I9525);
INV_X1 g_g5127 (I9525, g5127);
INV_X1 g_I9528 (g4006, I9528);
INV_X1 g_g5128 (I9528, g5128);
INV_X1 g_I9531 (g4463, I9531);
INV_X1 g_g5129 (I9531, g5129);
INV_X1 g_I9539 (g4018, I9539);
INV_X1 g_g5137 (I9539, g5137);
INV_X1 g_I9543 (g4279, I9543);
INV_X1 g_g5139 (I9543, g5139);
INV_X1 g_I9555 (g4892, I9555);
INV_X1 g_g5143 (I9555, g5143);
INV_X1 g_I9558 (g4597, I9558);
INV_X1 g_g5144 (I9558, g5144);
INV_X1 g_I9561 (g4695, I9561);
INV_X1 g_g5145 (I9561, g5145);
INV_X1 g_I9564 (g4703, I9564);
INV_X1 g_g5146 (I9564, g5146);
INV_X1 g_I9567 (g4693, I9567);
INV_X1 g_g5147 (I9567, g5147);
INV_X1 g_I9570 (g4696, I9570);
INV_X1 g_g5148 (I9570, g5148);
INV_X1 g_I9573 (g4701, I9573);
INV_X1 g_g5149 (I9573, g5149);
INV_X1 g_I9576 (g4706, I9576);
INV_X1 g_g5150 (I9576, g5150);
INV_X1 g_I9579 (g4713, I9579);
INV_X1 g_g5151 (I9579, g5151);
INV_X1 g_I9582 (g4694, I9582);
INV_X1 g_g5152 (I9582, g5152);
INV_X1 g_I9585 (g4697, I9585);
INV_X1 g_g5153 (I9585, g5153);
INV_X1 g_I9588 (g4704, I9588);
INV_X1 g_g5154 (I9588, g5154);
INV_X1 g_I9591 (g4710, I9591);
INV_X1 g_g5155 (I9591, g5155);
INV_X1 g_I9594 (g4718, I9594);
INV_X1 g_g5156 (I9594, g5156);
INV_X1 g_I9597 (g4738, I9597);
INV_X1 g_g5157 (I9597, g5157);
INV_X1 g_I9600 (g4698, I9600);
INV_X1 g_g5158 (I9600, g5158);
INV_X1 g_I9603 (g4719, I9603);
INV_X1 g_g5159 (I9603, g5159);
INV_X1 g_I9606 (g4687, I9606);
INV_X1 g_g5160 (I9606, g5160);
INV_X1 g_I9609 (g4780, I9609);
INV_X1 g_g5161 (I9609, g5161);
INV_X1 g_I9612 (g4776, I9612);
INV_X1 g_g5162 (I9612, g5162);
INV_X1 g_I9615 (g4739, I9615);
INV_X1 g_g5163 (I9615, g5163);
INV_X1 g_I9618 (g4742, I9618);
INV_X1 g_g5164 (I9618, g5164);
INV_X1 g_I9621 (g4732, I9621);
INV_X1 g_g5165 (I9621, g5165);
INV_X1 g_I9624 (g4746, I9624);
INV_X1 g_g5166 (I9624, g5166);
INV_X1 g_I9627 (g4777, I9627);
INV_X1 g_g5167 (I9627, g5167);
INV_X1 g_I9630 (g4867, I9630);
INV_X1 g_g5168 (I9630, g5168);
INV_X1 g_I9633 (g4800, I9633);
INV_X1 g_g5169 (I9633, g5169);
INV_X1 g_I9636 (g4802, I9636);
INV_X1 g_g5170 (I9636, g5170);
INV_X1 g_I9639 (g4685, I9639);
INV_X1 g_g5171 (I9639, g5171);
INV_X1 g_I9642 (g4788, I9642);
INV_X1 g_g5172 (I9642, g5172);
INV_X1 g_I9645 (g4900, I9645);
INV_X1 g_g5173 (I9645, g5173);
INV_X1 g_I9648 (g4795, I9648);
INV_X1 g_g5174 (I9648, g5174);
INV_X1 g_I9651 (g4805, I9651);
INV_X1 g_g5175 (I9651, g5175);
INV_X1 g_I9654 (g4792, I9654);
INV_X1 g_g5176 (I9654, g5176);
INV_X1 g_I9657 (g4784, I9657);
INV_X1 g_g5177 (I9657, g5177);
INV_X1 g_I9660 (g4806, I9660);
INV_X1 g_g5178 (I9660, g5178);
INV_X1 g_I9663 (g4809, I9663);
INV_X1 g_g5179 (I9663, g5179);
INV_X1 g_I9666 (g4931, I9666);
INV_X1 g_g5180 (I9666, g5180);
INV_X1 g_I9669 (g4909, I9669);
INV_X1 g_g5181 (I9669, g5181);
INV_X1 g_I9672 (g4803, I9672);
INV_X1 g_g5182 (I9672, g5182);
INV_X1 g_I9675 (g4807, I9675);
INV_X1 g_g5183 (I9675, g5183);
INV_X1 g_I9678 (g4808, I9678);
INV_X1 g_g5184 (I9678, g5184);
INV_X1 g_I9681 (g4811, I9681);
INV_X1 g_g5185 (I9681, g5185);
INV_X1 g_I9684 (g4813, I9684);
INV_X1 g_g5186 (I9684, g5186);
INV_X1 g_I9687 (g4822, I9687);
INV_X1 g_g5187 (I9687, g5187);
INV_X1 g_g5190 (g4938, g5190);
INV_X1 g_g5191 (g4969, g5191);
INV_X1 g_g5192 (g4841, g5192);
INV_X1 g_g5197 (g4938, g5197);
INV_X1 g_g5198 (g4969, g5198);
INV_X1 g_g5199 (g4841, g5199);
INV_X1 g_g5206 (g4938, g5206);
INV_X1 g_g5207 (g4673, g5207);
INV_X1 g_g5224 (g5114, g5224);
INV_X1 g_I9752 (g4705, I9752);
INV_X1 g_g5240 (I9752, g5240);
INV_X1 g_I9760 (g4838, I9760);
INV_X1 g_g5246 (I9760, g5246);
INV_X1 g_I9774 (g4678, I9774);
INV_X1 g_g5258 (I9774, g5258);
INV_X1 g_g5261 (g4748, g5261);
INV_X1 g_I9782 (g4720, I9782);
INV_X1 g_g5266 (I9782, g5266);
INV_X1 g_I9785 (g4747, I9785);
INV_X1 g_g5267 (I9785, g5267);
INV_X1 g_I9788 (g4711, I9788);
INV_X1 g_g5268 (I9788, g5268);
INV_X1 g_I9791 (g4779, I9791);
INV_X1 g_g5269 (I9791, g5269);
INV_X1 g_I9794 (g4778, I9794);
INV_X1 g_g5278 (I9794, g5278);
INV_X1 g_g5285 (g4841, g5285);
INV_X1 g_g5286 (g4714, g5286);
INV_X1 g_g5294 (g5087, g5294);
INV_X1 g_I9804 (g5113, I9804);
INV_X1 g_g5299 (I9804, g5299);
INV_X1 g_g5302 (g5028, g5302);
INV_X1 g_g5309 (g4969, g5309);
INV_X1 g_g5311 (g4938, g5311);
INV_X1 g_g5335 (g4677, g5335);
INV_X1 g_I9819 (g4691, I9819);
INV_X1 g_g5344 (I9819, g5344);
INV_X1 g_I9823 (g5138, I9823);
INV_X1 g_g5362 (I9823, g5362);
INV_X1 g_g5364 (g5124, g5364);
INV_X1 g_I9834 (g4782, I9834);
INV_X1 g_g5367 (I9834, g5367);
INV_X1 g_I9837 (g4781, I9837);
INV_X1 g_g5384 (I9837, g5384);
INV_X1 g_I9840 (g4702, I9840);
INV_X1 g_g5395 (I9840, g5395);
INV_X1 g_g5396 (g4692, g5396);
INV_X1 g_g5397 (g5076, g5397);
INV_X1 g_I9845 (g4728, I9845);
INV_X1 g_g5401 (I9845, g5401);
INV_X1 g_g5402 (g5000, g5402);
INV_X1 g_g5403 (g5088, g5403);
INV_X1 g_I9850 (g4798, I9850);
INV_X1 g_g5412 (I9850, g5412);
INV_X1 g_g5417 (g5006, g5417);
INV_X1 g_g5418 (g5100, g5418);
INV_X1 g_g5426 (g5013, g5426);
INV_X1 g_g5427 (g5115, g5427);
INV_X1 g_g5433 (g5024, g5433);
INV_X1 g_g5434 (g5112, g5434);
INV_X1 g_g5435 (g5121, g5435);
INV_X1 g_g5437 (g5041, g5437);
INV_X1 g_g5439 (g5058, g5439);
INV_X1 g_g5444 (g5074, g5444);
INV_X1 g_g5445 (g5059, g5445);
INV_X1 g_g5448 (g5137, g5448);
INV_X1 g_g5453 (g4680, g5453);
INV_X1 g_g5459 (g4882, g5459);
INV_X1 g_g5460 (g4684, g5460);
INV_X1 g_g5461 (g4885, g5461);
INV_X1 g_g5462 (g4886, g5462);
INV_X1 g_g5463 (g5085, g5463);
INV_X1 g_g5466 (g4890, g5466);
INV_X1 g_g5467 (g4891, g5467);
INV_X1 g_I9884 (g4868, I9884);
INV_X1 g_g5468 (I9884, g5468);
INV_X1 g_g5469 (g4898, g5469);
INV_X1 g_g5470 (g4899, g5470);
INV_X1 g_I9889 (g4819, I9889);
INV_X1 g_g5471 (I9889, g5471);
INV_X1 g_I9892 (g4879, I9892);
INV_X1 g_g5472 (I9892, g5472);
INV_X1 g_g5473 (g4903, g5473);
INV_X1 g_g5474 (g4904, g5474);
INV_X1 g_g5476 (g4907, g5476);
INV_X1 g_g5477 (g4908, g5477);
INV_X1 g_g5478 (g5025, g5478);
INV_X1 g_g5480 (g4913, g5480);
INV_X1 g_g5481 (g4914, g5481);
INV_X1 g_g5482 (g4915, g5482);
INV_X1 g_I9907 (g4837, I9907);
INV_X1 g_g5487 (I9907, g5487);
INV_X1 g_I9910 (g4681, I9910);
INV_X1 g_g5488 (I9910, g5488);
INV_X1 g_g5490 (g4917, g5490);
INV_X1 g_g5491 (g4918, g5491);
INV_X1 g_g5492 (g4919, g5492);
INV_X1 g_g5493 (g4920, g5493);
INV_X1 g_I9918 (g4968, I9918);
INV_X1 g_g5494 (I9918, g5494);
INV_X1 g_g5514 (g4922, g5514);
INV_X1 g_g5515 (g4923, g5515);
INV_X1 g_g5516 (g4924, g5516);
INV_X1 g_g5517 (g4925, g5517);
INV_X1 g_I9929 (g5052, I9929);
INV_X1 g_g5519 (I9929, g5519);
INV_X1 g_g5520 (g4928, g5520);
INV_X1 g_g5521 (g4929, g5521);
INV_X1 g_g5522 (g4930, g5522);
INV_X1 g_I9935 (g4812, I9935);
INV_X1 g_g5523 (I9935, g5523);
INV_X1 g_I9938 (g4878, I9938);
INV_X1 g_g5524 (I9938, g5524);
INV_X1 g_g5525 (g4934, g5525);
INV_X1 g_g5526 (g5086, g5526);
INV_X1 g_g5529 (g4689, g5529);
INV_X1 g_g5541 (g4814, g5541);
INV_X1 g_g5542 (g5061, g5542);
INV_X1 g_I9974 (g4676, I9974);
INV_X1 g_g5551 (I9974, g5551);
INV_X1 g_I10028 (g4825, I10028);
INV_X1 g_g5569 (I10028, g5569);
INV_X1 g_I10032 (g1236, I10032);
INV_X1 g_g5571 (I10032, g5571);
INV_X1 g_g5574 (g4969, g5574);
INV_X1 g_I10046 (g4840, I10046);
INV_X1 g_g5577 (I10046, g5577);
INV_X1 g_g5578 (g4841, g5578);
INV_X1 g_g5580 (g4938, g5580);
INV_X1 g_g5581 (g4969, g5581);
INV_X1 g_g5582 (g4969, g5582);
INV_X1 g_g5584 (g4841, g5584);
INV_X1 g_g5586 (g4938, g5586);
INV_X1 g_g5587 (g4938, g5587);
INV_X1 g_g5591 (g4841, g5591);
INV_X1 g_g5592 (g4969, g5592);
INV_X1 g_g5596 (g4841, g5596);
INV_X1 g_g5597 (g4969, g5597);
INV_X1 g_g5598 (g4938, g5598);
INV_X1 g_g5600 (g5128, g5600);
INV_X1 g_g5603 (g4938, g5603);
INV_X1 g_g5604 (g4969, g5604);
INV_X1 g_g5606 (g4748, g5606);
INV_X1 g_g5607 (g4938, g5607);
INV_X1 g_g5608 (g4969, g5608);
INV_X1 g_g5609 (g4748, g5609);
INV_X1 g_g5610 (g4938, g5610);
INV_X1 g_g5611 (g4969, g5611);
INV_X1 g_g5612 (g4814, g5612);
INV_X1 g_g5613 (g4748, g5613);
INV_X1 g_g5616 (g4938, g5616);
INV_X1 g_g5617 (g4969, g5617);
INV_X1 g_g5618 (g5015, g5618);
INV_X1 g_g5621 (g4748, g5621);
INV_X1 g_g5622 (g4938, g5622);
INV_X1 g_g5623 (g4969, g5623);
INV_X1 g_g5626 (g4748, g5626);
INV_X1 g_g5627 (g4673, g5627);
INV_X1 g_g5628 (g4748, g5628);
INV_X1 g_g5631 (g4938, g5631);
INV_X1 g_g5633 (g4895, g5633);
INV_X1 g_g5638 (g4748, g5638);
INV_X1 g_g5639 (g4748, g5639);
INV_X1 g_I10125 (g5127, I10125);
INV_X1 g_g5642 (I10125, g5642);
INV_X1 g_I10128 (g4688, I10128);
INV_X1 g_g5643 (I10128, g5643);
INV_X1 g_g5644 (g4748, g5644);
INV_X1 g_g5645 (g4748, g5645);
INV_X1 g_g5648 (g4748, g5648);
INV_X1 g_g5649 (g4748, g5649);
INV_X1 g_I10135 (g4960, I10135);
INV_X1 g_g5652 (I10135, g5652);
INV_X1 g_g5653 (g4748, g5653);
INV_X1 g_g5654 (g4748, g5654);
INV_X1 g_g5658 (g4748, g5658);
INV_X1 g_g5662 (g5027, g5662);
INV_X1 g_g5665 (g4748, g5665);
INV_X1 g_I10151 (g5007, I10151);
INV_X1 g_g5668 (I10151, g5668);
INV_X1 g_I10154 (g5109, I10154);
INV_X1 g_g5669 (I10154, g5669);
INV_X1 g_I10157 (g5109, I10157);
INV_X1 g_g5670 (I10157, g5670);
INV_X1 g_I10160 (g5139, I10160);
INV_X1 g_g5671 (I10160, g5671);
INV_X1 g_g5674 (g5042, g5674);
INV_X1 g_I10166 (g5016, I10166);
INV_X1 g_g5677 (I10166, g5677);
INV_X1 g_I10169 (g4873, I10169);
INV_X1 g_g5678 (I10169, g5678);
INV_X1 g_I10172 (g4873, I10172);
INV_X1 g_g5679 (I10172, g5679);
INV_X1 g_g5680 (g5101, g5680);
INV_X1 g_I10177 (g4721, I10177);
INV_X1 g_g5682 (I10177, g5682);
INV_X1 g_I10180 (g4721, I10180);
INV_X1 g_g5683 (I10180, g5683);
INV_X1 g_I10183 (g5129, I10183);
INV_X1 g_g5684 (I10183, g5684);
INV_X1 g_I10186 (g5129, I10186);
INV_X1 g_g5685 (I10186, g5685);
INV_X1 g_I10190 (g4670, I10190);
INV_X1 g_g5687 (I10190, g5687);
INV_X1 g_I10193 (g4670, I10193);
INV_X1 g_g5688 (I10193, g5688);
INV_X1 g_g5690 (g4748, g5690);
INV_X1 g_I10204 (g5060, I10204);
INV_X1 g_g5693 (I10204, g5693);
INV_X1 g_I10207 (g5075, I10207);
INV_X1 g_g5696 (I10207, g5696);
INV_X1 g_g5701 (g5120, g5701);
INV_X1 g_g5705 (g4841, g5705);
INV_X1 g_g5709 (g4841, g5709);
INV_X1 g_g5713 (g4841, g5713);
INV_X1 g_g5717 (g4969, g5717);
INV_X1 g_g5718 (g4841, g5718);
INV_X1 g_I10236 (g5014, I10236);
INV_X1 g_g5719 (I10236, g5719);
INV_X1 g_g5723 (g4938, g5723);
INV_X1 g_g5724 (g4969, g5724);
INV_X1 g_g5725 (g4841, g5725);
INV_X1 g_I10243 (g5026, I10243);
INV_X1 g_g5726 (I10243, g5726);
INV_X1 g_g5729 (g5144, g5729);
INV_X1 g_I10247 (g5266, I10247);
INV_X1 g_g5730 (I10247, g5730);
INV_X1 g_I10250 (g5268, I10250);
INV_X1 g_g5731 (I10250, g5731);
INV_X1 g_I10253 (g5240, I10253);
INV_X1 g_g5732 (I10253, g5732);
INV_X1 g_I10256 (g5401, I10256);
INV_X1 g_g5733 (I10256, g5733);
INV_X1 g_I10259 (g5362, I10259);
INV_X1 g_g5734 (I10259, g5734);
INV_X1 g_I10262 (g5551, I10262);
INV_X1 g_g5735 (I10262, g5735);
INV_X1 g_I10265 (g5468, I10265);
INV_X1 g_g5736 (I10265, g5736);
INV_X1 g_I10268 (g5471, I10268);
INV_X1 g_g5737 (I10268, g5737);
INV_X1 g_I10271 (g5487, I10271);
INV_X1 g_g5738 (I10271, g5738);
INV_X1 g_I10274 (g5524, I10274);
INV_X1 g_g5739 (I10274, g5739);
INV_X1 g_I10277 (g5472, I10277);
INV_X1 g_g5740 (I10277, g5740);
INV_X1 g_I10280 (g5488, I10280);
INV_X1 g_g5741 (I10280, g5741);
INV_X1 g_I10283 (g5643, I10283);
INV_X1 g_g5742 (I10283, g5742);
INV_X1 g_I10286 (g5519, I10286);
INV_X1 g_g5743 (I10286, g5743);
INV_X1 g_I10289 (g5569, I10289);
INV_X1 g_g5744 (I10289, g5744);
INV_X1 g_I10292 (g5577, I10292);
INV_X1 g_g5745 (I10292, g5745);
INV_X1 g_I10295 (g5523, I10295);
INV_X1 g_g5746 (I10295, g5746);
INV_X1 g_g5749 (g5207, g5749);
INV_X1 g_g5754 (g5403, g5754);
INV_X1 g_g5755 (g5494, g5755);
INV_X1 g_I10343 (g5704, I10343);
INV_X1 g_g5756 (I10343, g5756);
INV_X1 g_g5757 (g5261, g5757);
INV_X1 g_I10347 (g5706, I10347);
INV_X1 g_g5758 (I10347, g5758);
INV_X1 g_I10350 (g5707, I10350);
INV_X1 g_g5759 (I10350, g5759);
INV_X1 g_I10353 (g5710, I10353);
INV_X1 g_g5760 (I10353, g5760);
INV_X1 g_I10356 (g5711, I10356);
INV_X1 g_g5761 (I10356, g5761);
INV_X1 g_I10366 (g5715, I10366);
INV_X1 g_g5763 (I10366, g5763);
INV_X1 g_I10369 (g5716, I10369);
INV_X1 g_g5764 (I10369, g5764);
INV_X1 g_I10373 (g5722, I10373);
INV_X1 g_g5766 (I10373, g5766);
INV_X1 g_I10377 (g5188, I10377);
INV_X1 g_g5768 (I10377, g5768);
INV_X1 g_I10380 (g5448, I10380);
INV_X1 g_g5769 (I10380, g5769);
INV_X1 g_I10384 (g5193, I10384);
INV_X1 g_g5779 (I10384, g5779);
INV_X1 g_I10387 (g5194, I10387);
INV_X1 g_g5780 (I10387, g5780);
INV_X1 g_I10390 (g5195, I10390);
INV_X1 g_g5781 (I10390, g5781);
INV_X1 g_I10393 (g5196, I10393);
INV_X1 g_g5782 (I10393, g5782);
INV_X1 g_I10397 (g5200, I10397);
INV_X1 g_g5784 (I10397, g5784);
INV_X1 g_I10400 (g5201, I10400);
INV_X1 g_g5785 (I10400, g5785);
INV_X1 g_I10403 (g5202, I10403);
INV_X1 g_g5786 (I10403, g5786);
INV_X1 g_I10406 (g5203, I10406);
INV_X1 g_g5787 (I10406, g5787);
INV_X1 g_I10409 (g5204, I10409);
INV_X1 g_g5788 (I10409, g5788);
INV_X1 g_I10412 (g5205, I10412);
INV_X1 g_g5789 (I10412, g5789);
INV_X1 g_I10415 (g5397, I10415);
INV_X1 g_g5790 (I10415, g5790);
INV_X1 g_I10418 (g5453, I10418);
INV_X1 g_g5793 (I10418, g5793);
INV_X1 g_I10421 (g5208, I10421);
INV_X1 g_g5794 (I10421, g5794);
INV_X1 g_I10424 (g5209, I10424);
INV_X1 g_g5795 (I10424, g5795);
INV_X1 g_I10427 (g5210, I10427);
INV_X1 g_g5796 (I10427, g5796);
INV_X1 g_I10430 (g5211, I10430);
INV_X1 g_g5797 (I10430, g5797);
INV_X1 g_I10433 (g5212, I10433);
INV_X1 g_g5798 (I10433, g5798);
INV_X1 g_I10436 (g5213, I10436);
INV_X1 g_g5799 (I10436, g5799);
INV_X1 g_I10439 (g5214, I10439);
INV_X1 g_g5800 (I10439, g5800);
INV_X1 g_I10442 (g5215, I10442);
INV_X1 g_g5801 (I10442, g5801);
INV_X1 g_I10445 (g5418, I10445);
INV_X1 g_g5802 (I10445, g5802);
INV_X1 g_I10448 (g5335, I10448);
INV_X1 g_g5805 (I10448, g5805);
INV_X1 g_I10451 (g5216, I10451);
INV_X1 g_g5806 (I10451, g5806);
INV_X1 g_I10454 (g5217, I10454);
INV_X1 g_g5807 (I10454, g5807);
INV_X1 g_I10457 (g5218, I10457);
INV_X1 g_g5808 (I10457, g5808);
INV_X1 g_I10460 (g5219, I10460);
INV_X1 g_g5809 (I10460, g5809);
INV_X1 g_I10463 (g5220, I10463);
INV_X1 g_g5810 (I10463, g5810);
INV_X1 g_I10466 (g5221, I10466);
INV_X1 g_g5811 (I10466, g5811);
INV_X1 g_I10469 (g5222, I10469);
INV_X1 g_g5812 (I10469, g5812);
INV_X1 g_I10472 (g5223, I10472);
INV_X1 g_g5813 (I10472, g5813);
INV_X1 g_I10475 (g5529, I10475);
INV_X1 g_g5814 (I10475, g5814);
INV_X1 g_I10479 (g5227, I10479);
INV_X1 g_g5818 (I10479, g5818);
INV_X1 g_I10482 (g5228, I10482);
INV_X1 g_g5819 (I10482, g5819);
INV_X1 g_I10485 (g5229, I10485);
INV_X1 g_g5820 (I10485, g5820);
INV_X1 g_I10488 (g5230, I10488);
INV_X1 g_g5821 (I10488, g5821);
INV_X1 g_I10491 (g5231, I10491);
INV_X1 g_g5822 (I10491, g5822);
INV_X1 g_I10494 (g5232, I10494);
INV_X1 g_g5823 (I10494, g5823);
INV_X1 g_I10497 (g5233, I10497);
INV_X1 g_g5824 (I10497, g5824);
INV_X1 g_I10500 (g5234, I10500);
INV_X1 g_g5825 (I10500, g5825);
INV_X1 g_I10503 (g5235, I10503);
INV_X1 g_g5826 (I10503, g5826);
INV_X1 g_I10506 (g5236, I10506);
INV_X1 g_g5827 (I10506, g5827);
INV_X1 g_I10509 (g5237, I10509);
INV_X1 g_g5828 (I10509, g5828);
INV_X1 g_I10512 (g5238, I10512);
INV_X1 g_g5829 (I10512, g5829);
INV_X1 g_I10516 (g5241, I10516);
INV_X1 g_g5831 (I10516, g5831);
INV_X1 g_I10519 (g5242, I10519);
INV_X1 g_g5832 (I10519, g5832);
INV_X1 g_I10522 (g5243, I10522);
INV_X1 g_g5833 (I10522, g5833);
INV_X1 g_I10525 (g5244, I10525);
INV_X1 g_g5834 (I10525, g5834);
INV_X1 g_I10528 (g5245, I10528);
INV_X1 g_g5835 (I10528, g5835);
INV_X1 g_g5836 (g5529, g5836);
INV_X1 g_I10532 (g5253, I10532);
INV_X1 g_g5839 (I10532, g5839);
INV_X1 g_I10535 (g5254, I10535);
INV_X1 g_g5840 (I10535, g5840);
INV_X1 g_I10538 (g5255, I10538);
INV_X1 g_g5841 (I10538, g5841);
INV_X1 g_I10541 (g5256, I10541);
INV_X1 g_g5842 (I10541, g5842);
INV_X1 g_g5843 (g5367, g5843);
INV_X1 g_I10545 (g5259, I10545);
INV_X1 g_g5844 (I10545, g5844);
INV_X1 g_I10548 (g5260, I10548);
INV_X1 g_g5845 (I10548, g5845);
INV_X1 g_g5846 (g5367, g5846);
INV_X1 g_I10552 (g5396, I10552);
INV_X1 g_g5847 (I10552, g5847);
INV_X1 g_I10555 (g5529, I10555);
INV_X1 g_g5868 (I10555, g5868);
INV_X1 g_I10558 (g5264, I10558);
INV_X1 g_g5871 (I10558, g5871);
INV_X1 g_I10561 (g5265, I10561);
INV_X1 g_g5872 (I10561, g5872);
INV_X1 g_g5873 (g5367, g5873);
INV_X1 g_I10565 (g5402, I10565);
INV_X1 g_g5874 (I10565, g5874);
INV_X1 g_I10569 (g5417, I10569);
INV_X1 g_g5897 (I10569, g5897);
INV_X1 g_g5916 (g5384, g5916);
INV_X1 g_g5917 (g5412, g5917);
INV_X1 g_I10574 (g5426, I10574);
INV_X1 g_g5918 (I10574, g5918);
INV_X1 g_g5938 (g5412, g5938);
INV_X1 g_I10579 (g5433, I10579);
INV_X1 g_g5939 (I10579, g5939);
INV_X1 g_I10582 (g5437, I10582);
INV_X1 g_g5956 (I10582, g5956);
INV_X1 g_I10587 (g5439, I10587);
INV_X1 g_g5971 (I10587, g5971);
INV_X1 g_g5987 (g5294, g5987);
INV_X1 g_I10592 (g5444, I10592);
INV_X1 g_g5988 (I10592, g5988);
INV_X1 g_g6004 (g5494, g6004);
INV_X1 g_g6007 (g5494, g6007);
INV_X1 g_g6008 (g5367, g6008);
INV_X1 g_I10605 (g5440, I10605);
INV_X1 g_g6009 (I10605, g6009);
INV_X1 g_I10608 (g5701, I10608);
INV_X1 g_g6010 (I10608, g6010);
INV_X1 g_g6011 (g5494, g6011);
INV_X1 g_g6012 (g5367, g6012);
INV_X1 g_I10614 (g5302, I10614);
INV_X1 g_g6014 (I10614, g6014);
INV_X1 g_I10617 (g5677, I10617);
INV_X1 g_g6015 (I10617, g6015);
INV_X1 g_g6018 (g5494, g6018);
INV_X1 g_g6019 (g5367, g6019);
INV_X1 g_g6020 (g5367, g6020);
INV_X1 g_g6024 (g5494, g6024);
INV_X1 g_g6025 (g5367, g6025);
INV_X1 g_g6026 (g5384, g6026);
INV_X1 g_g6027 (g5384, g6027);
INV_X1 g_g6028 (g5529, g6028);
INV_X1 g_g6032 (g5494, g6032);
INV_X1 g_g6033 (g5384, g6033);
INV_X1 g_I10639 (g5224, I10639);
INV_X1 g_g6034 (I10639, g6034);
INV_X1 g_g6035 (g5494, g6035);
INV_X1 g_I10643 (g5267, I10643);
INV_X1 g_g6036 (I10643, g6036);
INV_X1 g_I10646 (g5364, I10646);
INV_X1 g_g6037 (I10646, g6037);
INV_X1 g_I10649 (g5657, I10649);
INV_X1 g_g6038 (I10649, g6038);
INV_X1 g_g6048 (g5246, g6048);
INV_X1 g_g6050 (g5246, g6050);
INV_X1 g_g6051 (g5246, g6051);
INV_X1 g_g6059 (g5317, g6059);
INV_X1 g_I10675 (g5662, I10675);
INV_X1 g_g6062 (I10675, g6062);
INV_X1 g_I10678 (g5566, I10678);
INV_X1 g_g6063 (I10678, g6063);
INV_X1 g_I10681 (g5686, I10681);
INV_X1 g_g6064 (I10681, g6064);
INV_X1 g_I10684 (g5258, I10684);
INV_X1 g_g6065 (I10684, g6065);
INV_X1 g_I10687 (g5674, I10687);
INV_X1 g_g6068 (I10687, g6068);
INV_X1 g_I10690 (g5538, I10690);
INV_X1 g_g6069 (I10690, g6069);
INV_X1 g_g6070 (g5317, g6070);
INV_X1 g_I10694 (g5445, I10694);
INV_X1 g_g6071 (I10694, g6071);
INV_X1 g_g6072 (g5345, g6072);
INV_X1 g_g6073 (g5384, g6073);
INV_X1 g_g6074 (g5317, g6074);
INV_X1 g_g6075 (g5345, g6075);
INV_X1 g_g6076 (g5287, g6076);
INV_X1 g_I10702 (g5529, I10702);
INV_X1 g_g6083 (I10702, g6083);
INV_X1 g_I10705 (g5463, I10705);
INV_X1 g_g6087 (I10705, g6087);
INV_X1 g_I10708 (g5545, I10708);
INV_X1 g_g6088 (I10708, g6088);
INV_X1 g_g6089 (g5317, g6089);
INV_X1 g_g6090 (g5529, g6090);
INV_X1 g_g6092 (g5317, g6092);
INV_X1 g_g6093 (g5345, g6093);
INV_X1 g_I10716 (g5537, I10716);
INV_X1 g_g6094 (I10716, g6094);
INV_X1 g_I10719 (g5559, I10719);
INV_X1 g_g6095 (I10719, g6095);
INV_X1 g_g6096 (g5317, g6096);
INV_X1 g_g6097 (g5345, g6097);
INV_X1 g_g6101 (g5317, g6101);
INV_X1 g_g6102 (g5345, g6102);
INV_X1 g_g6103 (g5317, g6103);
INV_X1 g_g6104 (g5345, g6104);
INV_X1 g_g6106 (g5345, g6106);
INV_X1 g_g6108 (g5345, g6108);
INV_X1 g_g6110 (g5335, g6110);
INV_X1 g_g6111 (g5453, g6111);
INV_X1 g_I10739 (g5572, I10739);
INV_X1 g_g6117 (I10739, g6117);
INV_X1 g_g6118 (g5549, g6118);
INV_X1 g_I10752 (g5618, I10752);
INV_X1 g_g6122 (I10752, g6122);
INV_X1 g_I10758 (g5662, I10758);
INV_X1 g_g6129 (I10758, g6129);
INV_X1 g_I10761 (g5302, I10761);
INV_X1 g_g6130 (I10761, g6130);
INV_X1 g_g6131 (g5529, g6131);
INV_X1 g_I10766 (g5674, I10766);
INV_X1 g_g6133 (I10766, g6133);
INV_X1 g_g6134 (g5428, g6134);
INV_X1 g_I10770 (g5441, I10770);
INV_X1 g_g6135 (I10770, g6135);
INV_X1 g_I10773 (g5708, I10773);
INV_X1 g_g6136 (I10773, g6136);
INV_X1 g_I10776 (g5576, I10776);
INV_X1 g_g6137 (I10776, g6137);
INV_X1 g_I10780 (g5445, I10780);
INV_X1 g_g6139 (I10780, g6139);
INV_X1 g_I10783 (g5542, I10783);
INV_X1 g_g6140 (I10783, g6140);
INV_X1 g_I10786 (g5452, I10786);
INV_X1 g_g6141 (I10786, g6141);
INV_X1 g_I10796 (g5397, I10796);
INV_X1 g_g6143 (I10796, g6143);
INV_X1 g_I10801 (g5463, I10801);
INV_X1 g_g6146 (I10801, g6146);
INV_X1 g_I10804 (g5526, I10804);
INV_X1 g_g6147 (I10804, g6147);
INV_X1 g_I10807 (g5294, I10807);
INV_X1 g_g6148 (I10807, g6148);
INV_X1 g_I10810 (g5403, I10810);
INV_X1 g_g6149 (I10810, g6149);
INV_X1 g_g6150 (g5287, g6150);
INV_X1 g_I10815 (g5418, I10815);
INV_X1 g_g6152 (I10815, g6152);
INV_X1 g_I10826 (g5434, I10826);
INV_X1 g_g6155 (I10826, g6155);
INV_X1 g_I10829 (g5224, I10829);
INV_X1 g_g6156 (I10829, g6156);
INV_X1 g_I10842 (g5701, I10842);
INV_X1 g_g6161 (I10842, g6161);
INV_X1 g_I10862 (g5364, I10862);
INV_X1 g_g6167 (I10862, g6167);
INV_X1 g_I10882 (g5600, I10882);
INV_X1 g_g6173 (I10882, g6173);
INV_X1 g_I10896 (g5475, I10896);
INV_X1 g_g6179 (I10896, g6179);
INV_X1 g_I10914 (g5448, I10914);
INV_X1 g_g6183 (I10914, g6183);
INV_X1 g_I10919 (g5479, I10919);
INV_X1 g_g6186 (I10919, g6186);
INV_X1 g_I10930 (g5600, I10930);
INV_X1 g_g6189 (I10930, g6189);
INV_X1 g_I10933 (g5668, I10933);
INV_X1 g_g6190 (I10933, g6190);
INV_X1 g_I10937 (g5560, I10937);
INV_X1 g_g6194 (I10937, g6194);
INV_X1 g_I10940 (g5489, I10940);
INV_X1 g_g6195 (I10940, g6195);
INV_X1 g_g6198 (g5335, g6198);
INV_X1 g_I10946 (g5563, I10946);
INV_X1 g_g6201 (I10946, g6201);
INV_X1 g_I10949 (g5513, I10949);
INV_X1 g_g6202 (I10949, g6202);
INV_X1 g_g6205 (g5628, g6205);
INV_X1 g_g6206 (g5639, g6206);
INV_X1 g_I10962 (g5719, I10962);
INV_X1 g_g6207 (I10962, g6207);
INV_X1 g_I10965 (g5719, I10965);
INV_X1 g_g6208 (I10965, g6208);
INV_X1 g_I10969 (g5606, I10969);
INV_X1 g_g6210 (I10969, g6210);
INV_X1 g_g6211 (g5645, g6211);
INV_X1 g_I10973 (g5726, I10973);
INV_X1 g_g6212 (I10973, g6212);
INV_X1 g_I10976 (g5726, I10976);
INV_X1 g_g6213 (I10976, g6213);
INV_X1 g_I10987 (g5609, I10987);
INV_X1 g_g6216 (I10987, g6216);
INV_X1 g_g6217 (g5649, g6217);
INV_X1 g_I10998 (g5672, I10998);
INV_X1 g_g6219 (I10998, g6219);
INV_X1 g_I11001 (g5698, I11001);
INV_X1 g_g6220 (I11001, g6220);
INV_X1 g_I11004 (g5613, I11004);
INV_X1 g_g6221 (I11004, g6221);
INV_X1 g_g6222 (g5654, g6222);
INV_X1 g_I11008 (g5693, I11008);
INV_X1 g_g6223 (I11008, g6223);
INV_X1 g_I11011 (g5693, I11011);
INV_X1 g_g6224 (I11011, g6224);
INV_X1 g_I11014 (g5621, I11014);
INV_X1 g_g6225 (I11014, g6225);
INV_X1 g_g6226 (g5658, g6226);
INV_X1 g_I11018 (g5626, I11018);
INV_X1 g_g6227 (I11018, g6227);
INV_X1 g_I11021 (g5627, I11021);
INV_X1 g_g6228 (I11021, g6228);
INV_X1 g_g6229 (g5665, g6229);
INV_X1 g_I11025 (g5638, I11025);
INV_X1 g_g6230 (I11025, g6230);
INV_X1 g_I11028 (g5642, I11028);
INV_X1 g_g6231 (I11028, g6231);
INV_X1 g_I11031 (g5335, I11031);
INV_X1 g_g6232 (I11031, g6232);
INV_X1 g_I11034 (g5644, I11034);
INV_X1 g_g6235 (I11034, g6235);
INV_X1 g_I11037 (g5299, I11037);
INV_X1 g_g6236 (I11037, g6236);
INV_X1 g_I11040 (g5299, I11040);
INV_X1 g_g6237 (I11040, g6237);
INV_X1 g_I11043 (g5648, I11043);
INV_X1 g_g6238 (I11043, g6238);
INV_X1 g_I11047 (g5653, I11047);
INV_X1 g_g6242 (I11047, g6242);
INV_X1 g_I11050 (g5335, I11050);
INV_X1 g_g6243 (I11050, g6243);
INV_X1 g_g6244 (g5670, g6244);
INV_X1 g_g6245 (g5690, g6245);
INV_X1 g_I11055 (g5696, I11055);
INV_X1 g_g6246 (I11055, g6246);
INV_X1 g_g6250 (g5679, g6250);
INV_X1 g_I11060 (g5453, I11060);
INV_X1 g_g6251 (I11060, g6251);
INV_X1 g_g6252 (g5418, g6252);
INV_X1 g_g6253 (g5403, g6253);
INV_X1 g_g6254 (g5683, g6254);
INV_X1 g_I11066 (g5460, I11066);
INV_X1 g_g6255 (I11066, g6255);
INV_X1 g_I11069 (g5671, I11069);
INV_X1 g_g6256 (I11069, g6256);
INV_X1 g_g6257 (g5685, g6257);
INV_X1 g_g6258 (g5427, g6258);
INV_X1 g_g6263 (g5688, g6263);
INV_X1 g_g6264 (g5403, g6264);
INV_X1 g_I11086 (g5397, I11086);
INV_X1 g_g6267 (I11086, g6267);
INV_X1 g_I11090 (g1000, I11090);
INV_X1 g_g6269 (I11090, g6269);
INV_X1 g_I11129 (g5418, I11129);
INV_X1 g_g6278 (I11129, g6278);
INV_X1 g_I11132 (g5624, I11132);
INV_X1 g_g6279 (I11132, g6279);
INV_X1 g_I11191 (g6155, I11191);
INV_X1 g_g6288 (I11191, g6288);
INV_X1 g_I11194 (g6243, I11194);
INV_X1 g_g6289 (I11194, g6289);
INV_X1 g_I11197 (g6122, I11197);
INV_X1 g_g6290 (I11197, g6290);
INV_X1 g_I11200 (g6251, I11200);
INV_X1 g_g6291 (I11200, g6291);
INV_X1 g_I11203 (g6129, I11203);
INV_X1 g_g6292 (I11203, g6292);
INV_X1 g_I11206 (g6133, I11206);
INV_X1 g_g6293 (I11206, g6293);
INV_X1 g_I11209 (g6139, I11209);
INV_X1 g_g6294 (I11209, g6294);
INV_X1 g_I11212 (g6146, I11212);
INV_X1 g_g6295 (I11212, g6295);
INV_X1 g_I11215 (g6156, I11215);
INV_X1 g_g6296 (I11215, g6296);
INV_X1 g_I11218 (g6161, I11218);
INV_X1 g_g6297 (I11218, g6297);
INV_X1 g_I11221 (g6167, I11221);
INV_X1 g_g6298 (I11221, g6298);
INV_X1 g_I11224 (g6255, I11224);
INV_X1 g_g6299 (I11224, g6299);
INV_X1 g_I11227 (g6130, I11227);
INV_X1 g_g6300 (I11227, g6300);
INV_X1 g_I11230 (g6140, I11230);
INV_X1 g_g6301 (I11230, g6301);
INV_X1 g_I11233 (g6147, I11233);
INV_X1 g_g6302 (I11233, g6302);
INV_X1 g_I11236 (g6148, I11236);
INV_X1 g_g6303 (I11236, g6303);
INV_X1 g_I11239 (g6173, I11239);
INV_X1 g_g6304 (I11239, g6304);
INV_X1 g_I11242 (g6183, I11242);
INV_X1 g_g6305 (I11242, g6305);
INV_X1 g_I11245 (g6143, I11245);
INV_X1 g_g6306 (I11245, g6306);
INV_X1 g_I11248 (g6149, I11248);
INV_X1 g_g6307 (I11248, g6307);
INV_X1 g_I11251 (g6152, I11251);
INV_X1 g_g6308 (I11251, g6308);
INV_X1 g_I11254 (g5793, I11254);
INV_X1 g_g6309 (I11254, g6309);
INV_X1 g_I11257 (g5805, I11257);
INV_X1 g_g6310 (I11257, g6310);
INV_X1 g_I11260 (g5779, I11260);
INV_X1 g_g6311 (I11260, g6311);
INV_X1 g_I11263 (g5784, I11263);
INV_X1 g_g6312 (I11263, g6312);
INV_X1 g_I11266 (g5794, I11266);
INV_X1 g_g6313 (I11266, g6313);
INV_X1 g_I11269 (g5756, I11269);
INV_X1 g_g6314 (I11269, g6314);
INV_X1 g_I11272 (g5758, I11272);
INV_X1 g_g6315 (I11272, g6315);
INV_X1 g_I11275 (g5768, I11275);
INV_X1 g_g6316 (I11275, g6316);
INV_X1 g_I11278 (g5780, I11278);
INV_X1 g_g6317 (I11278, g6317);
INV_X1 g_I11281 (g5785, I11281);
INV_X1 g_g6318 (I11281, g6318);
INV_X1 g_I11284 (g5795, I11284);
INV_X1 g_g6319 (I11284, g6319);
INV_X1 g_I11287 (g5806, I11287);
INV_X1 g_g6320 (I11287, g6320);
INV_X1 g_I11290 (g5818, I11290);
INV_X1 g_g6321 (I11290, g6321);
INV_X1 g_I11293 (g5824, I11293);
INV_X1 g_g6322 (I11293, g6322);
INV_X1 g_I11296 (g5831, I11296);
INV_X1 g_g6323 (I11296, g6323);
INV_X1 g_I11299 (g5786, I11299);
INV_X1 g_g6324 (I11299, g6324);
INV_X1 g_I11302 (g5796, I11302);
INV_X1 g_g6325 (I11302, g6325);
INV_X1 g_I11305 (g5807, I11305);
INV_X1 g_g6326 (I11305, g6326);
INV_X1 g_I11308 (g5759, I11308);
INV_X1 g_g6327 (I11308, g6327);
INV_X1 g_I11311 (g5760, I11311);
INV_X1 g_g6328 (I11311, g6328);
INV_X1 g_I11314 (g5781, I11314);
INV_X1 g_g6329 (I11314, g6329);
INV_X1 g_I11317 (g5787, I11317);
INV_X1 g_g6330 (I11317, g6330);
INV_X1 g_I11320 (g5797, I11320);
INV_X1 g_g6331 (I11320, g6331);
INV_X1 g_I11323 (g5808, I11323);
INV_X1 g_g6332 (I11323, g6332);
INV_X1 g_I11326 (g5819, I11326);
INV_X1 g_g6333 (I11326, g6333);
INV_X1 g_I11329 (g5825, I11329);
INV_X1 g_g6334 (I11329, g6334);
INV_X1 g_I11332 (g5832, I11332);
INV_X1 g_g6335 (I11332, g6335);
INV_X1 g_I11335 (g5839, I11335);
INV_X1 g_g6336 (I11335, g6336);
INV_X1 g_I11338 (g5798, I11338);
INV_X1 g_g6337 (I11338, g6337);
INV_X1 g_I11341 (g5809, I11341);
INV_X1 g_g6338 (I11341, g6338);
INV_X1 g_I11344 (g5820, I11344);
INV_X1 g_g6339 (I11344, g6339);
INV_X1 g_I11347 (g5761, I11347);
INV_X1 g_g6340 (I11347, g6340);
INV_X1 g_I11350 (g5763, I11350);
INV_X1 g_g6341 (I11350, g6341);
INV_X1 g_I11353 (g5788, I11353);
INV_X1 g_g6342 (I11353, g6342);
INV_X1 g_I11356 (g5799, I11356);
INV_X1 g_g6343 (I11356, g6343);
INV_X1 g_I11359 (g5810, I11359);
INV_X1 g_g6344 (I11359, g6344);
INV_X1 g_I11362 (g5821, I11362);
INV_X1 g_g6345 (I11362, g6345);
INV_X1 g_I11365 (g5826, I11365);
INV_X1 g_g6346 (I11365, g6346);
INV_X1 g_I11368 (g5833, I11368);
INV_X1 g_g6347 (I11368, g6347);
INV_X1 g_I11371 (g5840, I11371);
INV_X1 g_g6348 (I11371, g6348);
INV_X1 g_I11374 (g5844, I11374);
INV_X1 g_g6349 (I11374, g6349);
INV_X1 g_I11377 (g5811, I11377);
INV_X1 g_g6350 (I11377, g6350);
INV_X1 g_I11380 (g5822, I11380);
INV_X1 g_g6351 (I11380, g6351);
INV_X1 g_I11383 (g5827, I11383);
INV_X1 g_g6352 (I11383, g6352);
INV_X1 g_I11386 (g5764, I11386);
INV_X1 g_g6353 (I11386, g6353);
INV_X1 g_I11389 (g5766, I11389);
INV_X1 g_g6354 (I11389, g6354);
INV_X1 g_I11392 (g5800, I11392);
INV_X1 g_g6355 (I11392, g6355);
INV_X1 g_I11395 (g5812, I11395);
INV_X1 g_g6356 (I11395, g6356);
INV_X1 g_I11398 (g5823, I11398);
INV_X1 g_g6357 (I11398, g6357);
INV_X1 g_I11401 (g5828, I11401);
INV_X1 g_g6358 (I11401, g6358);
INV_X1 g_I11404 (g5834, I11404);
INV_X1 g_g6359 (I11404, g6359);
INV_X1 g_I11407 (g5841, I11407);
INV_X1 g_g6360 (I11407, g6360);
INV_X1 g_I11410 (g5845, I11410);
INV_X1 g_g6361 (I11410, g6361);
INV_X1 g_I11413 (g5871, I11413);
INV_X1 g_g6362 (I11413, g6362);
INV_X1 g_I11416 (g5829, I11416);
INV_X1 g_g6363 (I11416, g6363);
INV_X1 g_I11419 (g5835, I11419);
INV_X1 g_g6364 (I11419, g6364);
INV_X1 g_I11422 (g5842, I11422);
INV_X1 g_g6365 (I11422, g6365);
INV_X1 g_I11425 (g5872, I11425);
INV_X1 g_g6366 (I11425, g6366);
INV_X1 g_I11428 (g5813, I11428);
INV_X1 g_g6367 (I11428, g6367);
INV_X1 g_I11431 (g5782, I11431);
INV_X1 g_g6368 (I11431, g6368);
INV_X1 g_I11434 (g5789, I11434);
INV_X1 g_g6369 (I11434, g6369);
INV_X1 g_I11437 (g5801, I11437);
INV_X1 g_g6370 (I11437, g6370);
INV_X1 g_I11440 (g6009, I11440);
INV_X1 g_g6371 (I11440, g6371);
INV_X1 g_I11443 (g6038, I11443);
INV_X1 g_g6372 (I11443, g6372);
INV_X1 g_I11446 (g6062, I11446);
INV_X1 g_g6373 (I11446, g6373);
INV_X1 g_I11449 (g6068, I11449);
INV_X1 g_g6374 (I11449, g6374);
INV_X1 g_I11452 (g6071, I11452);
INV_X1 g_g6375 (I11452, g6375);
INV_X1 g_I11455 (g6087, I11455);
INV_X1 g_g6376 (I11455, g6376);
INV_X1 g_I11458 (g6063, I11458);
INV_X1 g_g6377 (I11458, g6377);
INV_X1 g_I11461 (g6094, I11461);
INV_X1 g_g6378 (I11461, g6378);
INV_X1 g_I11464 (g6088, I11464);
INV_X1 g_g6379 (I11464, g6379);
INV_X1 g_I11467 (g6064, I11467);
INV_X1 g_g6380 (I11467, g6380);
INV_X1 g_I11470 (g6095, I11470);
INV_X1 g_g6381 (I11470, g6381);
INV_X1 g_I11473 (g6069, I11473);
INV_X1 g_g6382 (I11473, g6382);
INV_X1 g_I11476 (g6194, I11476);
INV_X1 g_g6383 (I11476, g6383);
INV_X1 g_I11479 (g6201, I11479);
INV_X1 g_g6384 (I11479, g6384);
INV_X1 g_I11482 (g6117, I11482);
INV_X1 g_g6385 (I11482, g6385);
INV_X1 g_I11485 (g6137, I11485);
INV_X1 g_g6386 (I11485, g6386);
INV_X1 g_I11488 (g6034, I11488);
INV_X1 g_g6387 (I11488, g6387);
INV_X1 g_I11491 (g6010, I11491);
INV_X1 g_g6388 (I11491, g6388);
INV_X1 g_I11494 (g6037, I11494);
INV_X1 g_g6389 (I11494, g6389);
INV_X1 g_I11497 (g6014, I11497);
INV_X1 g_g6390 (I11497, g6390);
INV_X1 g_I11500 (g6219, I11500);
INV_X1 g_g6391 (I11500, g6391);
INV_X1 g_I11503 (g6220, I11503);
INV_X1 g_g6392 (I11503, g6392);
INV_X1 g_I11506 (g6189, I11506);
INV_X1 g_g6393 (I11506, g6393);
INV_X1 g_I11512 (g5874, I11512);
INV_X1 g_g6397 (I11512, g6397);
INV_X1 g_I11515 (g5897, I11515);
INV_X1 g_g6398 (I11515, g6398);
INV_X1 g_I11522 (g5847, I11522);
INV_X1 g_g6403 (I11522, g6403);
INV_X1 g_I11525 (g5874, I11525);
INV_X1 g_g6404 (I11525, g6404);
INV_X1 g_I11533 (g5847, I11533);
INV_X1 g_g6410 (I11533, g6410);
INV_X1 g_I11556 (g6065, I11556);
INV_X1 g_g6425 (I11556, g6425);
INV_X1 g_I11559 (g6065, I11559);
INV_X1 g_g6426 (I11559, g6426);
INV_X1 g_I11562 (g5939, I11562);
INV_X1 g_g6427 (I11562, g6427);
INV_X1 g_I11569 (g6279, I11569);
INV_X1 g_g6432 (I11569, g6432);
INV_X1 g_I11586 (g6256, I11586);
INV_X1 g_g6441 (I11586, g6441);
INV_X1 g_I11591 (g5814, I11591);
INV_X1 g_g6446 (I11591, g6446);
INV_X1 g_I11596 (g6228, I11596);
INV_X1 g_g6449 (I11596, g6449);
INV_X1 g_I11607 (g5767, I11607);
INV_X1 g_g6461 (I11607, g6461);
INV_X1 g_I11622 (g5847, I11622);
INV_X1 g_g6468 (I11622, g6468);
INV_X1 g_I11627 (g5874, I11627);
INV_X1 g_g6471 (I11627, g6471);
INV_X1 g_I11633 (g5897, I11633);
INV_X1 g_g6475 (I11633, g6475);
INV_X1 g_I11638 (g5847, I11638);
INV_X1 g_g6478 (I11638, g6478);
INV_X1 g_I11641 (g5918, I11641);
INV_X1 g_g6481 (I11641, g6481);
INV_X1 g_I11645 (g5874, I11645);
INV_X1 g_g6483 (I11645, g6483);
INV_X1 g_I11648 (g6028, I11648);
INV_X1 g_g6486 (I11648, g6486);
INV_X1 g_I11652 (g5939, I11652);
INV_X1 g_g6488 (I11652, g6488);
INV_X1 g_I11656 (g5772, I11656);
INV_X1 g_g6490 (I11656, g6490);
INV_X1 g_I11659 (g5897, I11659);
INV_X1 g_g6493 (I11659, g6493);
INV_X1 g_I11662 (g5956, I11662);
INV_X1 g_g6496 (I11662, g6496);
INV_X1 g_I11666 (g5772, I11666);
INV_X1 g_g6498 (I11666, g6498);
INV_X1 g_I11669 (g5918, I11669);
INV_X1 g_g6501 (I11669, g6501);
INV_X1 g_I11672 (g5971, I11672);
INV_X1 g_g6502 (I11672, g6502);
INV_X1 g_I11677 (g6076, I11677);
INV_X1 g_g6505 (I11677, g6505);
INV_X1 g_I11680 (g5939, I11680);
INV_X1 g_g6506 (I11680, g6506);
INV_X1 g_I11683 (g5988, I11683);
INV_X1 g_g6507 (I11683, g6507);
INV_X1 g_I11686 (g6076, I11686);
INV_X1 g_g6508 (I11686, g6508);
INV_X1 g_I11689 (g5956, I11689);
INV_X1 g_g6509 (I11689, g6509);
INV_X1 g_I11693 (g6076, I11693);
INV_X1 g_g6511 (I11693, g6511);
INV_X1 g_I11696 (g5971, I11696);
INV_X1 g_g6514 (I11696, g6514);
INV_X1 g_g6515 (g6125, g6515);
INV_X1 g_I11701 (g5772, I11701);
INV_X1 g_g6517 (I11701, g6517);
INV_X1 g_I11704 (g6076, I11704);
INV_X1 g_g6520 (I11704, g6520);
INV_X1 g_I11707 (g5988, I11707);
INV_X1 g_g6523 (I11707, g6523);
INV_X1 g_I11710 (g6098, I11710);
INV_X1 g_g6524 (I11710, g6524);
INV_X1 g_I11714 (g5772, I11714);
INV_X1 g_g6538 (I11714, g6538);
INV_X1 g_I11718 (g6115, I11718);
INV_X1 g_g6542 (I11718, g6542);
INV_X1 g_I11722 (g5772, I11722);
INV_X1 g_g6552 (I11722, g6552);
INV_X1 g_I11725 (g6036, I11725);
INV_X1 g_g6553 (I11725, g6553);
INV_X1 g_I11729 (g5772, I11729);
INV_X1 g_g6555 (I11729, g6555);
INV_X1 g_I11732 (g6076, I11732);
INV_X1 g_g6556 (I11732, g6556);
INV_X1 g_I11736 (g6076, I11736);
INV_X1 g_g6562 (I11736, g6562);
INV_X1 g_I11740 (g6136, I11740);
INV_X1 g_g6566 (I11740, g6566);
INV_X1 g_I11744 (g6120, I11744);
INV_X1 g_g6568 (I11744, g6568);
INV_X1 g_I11747 (g6123, I11747);
INV_X1 g_g6569 (I11747, g6569);
INV_X1 g_I11764 (g6056, I11764);
INV_X1 g_g6572 (I11764, g6572);
INV_X1 g_g6573 (g5868, g6573);
INV_X1 g_I11773 (g6262, I11773);
INV_X1 g_g6581 (I11773, g6581);
INV_X1 g_I11778 (g6180, I11778);
INV_X1 g_g6586 (I11778, g6586);
INV_X1 g_I11781 (g6284, I11781);
INV_X1 g_g6587 (I11781, g6587);
INV_X1 g_g6588 (g5836, g6588);
INV_X1 g_g6589 (g6083, g6589);
INV_X1 g_I11787 (g6273, I11787);
INV_X1 g_g6591 (I11787, g6591);
INV_X1 g_I11790 (g6282, I11790);
INV_X1 g_g6592 (I11790, g6592);
INV_X1 g_I11793 (g6188, I11793);
INV_X1 g_g6593 (I11793, g6593);
INV_X1 g_I11796 (g6287, I11796);
INV_X1 g_g6594 (I11796, g6594);
INV_X1 g_g6595 (g6083, g6595);
INV_X1 g_I11800 (g6164, I11800);
INV_X1 g_g6596 (I11800, g6596);
INV_X1 g_I11803 (g6280, I11803);
INV_X1 g_g6597 (I11803, g6597);
INV_X1 g_I11806 (g6275, I11806);
INV_X1 g_g6598 (I11806, g6598);
INV_X1 g_I11809 (g6285, I11809);
INV_X1 g_g6599 (I11809, g6599);
INV_X1 g_g6601 (g6083, g6601);
INV_X1 g_I11815 (g6169, I11815);
INV_X1 g_g6603 (I11815, g6603);
INV_X1 g_I11818 (g6276, I11818);
INV_X1 g_g6604 (I11818, g6604);
INV_X1 g_I11821 (g6170, I11821);
INV_X1 g_g6605 (I11821, g6605);
INV_X1 g_I11824 (g6283, I11824);
INV_X1 g_g6606 (I11824, g6606);
INV_X1 g_I11827 (g6231, I11827);
INV_X1 g_g6607 (I11827, g6607);
INV_X1 g_I11832 (g6274, I11832);
INV_X1 g_g6612 (I11832, g6612);
INV_X1 g_I11835 (g6181, I11835);
INV_X1 g_g6613 (I11835, g6613);
INV_X1 g_I11838 (g6281, I11838);
INV_X1 g_g6614 (I11838, g6614);
INV_X1 g_I11848 (g6159, I11848);
INV_X1 g_g6616 (I11848, g6616);
INV_X1 g_I11851 (g6277, I11851);
INV_X1 g_g6617 (I11851, g6617);
INV_X1 g_g6618 (g6003, g6618);
INV_X1 g_I11855 (g5751, I11855);
INV_X1 g_g6621 (I11855, g6621);
INV_X1 g_I11858 (g6165, I11858);
INV_X1 g_g6622 (I11858, g6622);
INV_X1 g_I11861 (g5747, I11861);
INV_X1 g_g6623 (I11861, g6623);
INV_X1 g_I11864 (g5753, I11864);
INV_X1 g_g6624 (I11864, g6624);
INV_X1 g_I11867 (g6286, I11867);
INV_X1 g_g6625 (I11867, g6625);
INV_X1 g_I11870 (g5752, I11870);
INV_X1 g_g6626 (I11870, g6626);
INV_X1 g_I11880 (g5748, I11880);
INV_X1 g_g6628 (I11880, g6628);
INV_X1 g_I11884 (g6091, I11884);
INV_X1 g_g6630 (I11884, g6630);
INV_X1 g_I11887 (g5918, I11887);
INV_X1 g_g6631 (I11887, g6631);
INV_X1 g_I11890 (g6135, I11890);
INV_X1 g_g6632 (I11890, g6632);
INV_X1 g_I11894 (g5956, I11894);
INV_X1 g_g6634 (I11894, g6634);
INV_X1 g_I11897 (g6141, I11897);
INV_X1 g_g6635 (I11897, g6635);
INV_X1 g_I11900 (g5847, I11900);
INV_X1 g_g6636 (I11900, g6636);
INV_X1 g_I11903 (g5939, I11903);
INV_X1 g_g6637 (I11903, g6637);
INV_X1 g_g6639 (g6198, g6639);
INV_X1 g_I11908 (g5918, I11908);
INV_X1 g_g6640 (I11908, g6640);
INV_X1 g_I11912 (g5897, I11912);
INV_X1 g_g6642 (I11912, g6642);
INV_X1 g_g6644 (g6208, g6644);
INV_X1 g_I11917 (g5897, I11917);
INV_X1 g_g6645 (I11917, g6645);
INV_X1 g_I11920 (g5874, I11920);
INV_X1 g_g6646 (I11920, g6646);
INV_X1 g_I11923 (g5939, I11923);
INV_X1 g_g6647 (I11923, g6647);
INV_X1 g_I11926 (g6190, I11926);
INV_X1 g_g6648 (I11926, g6648);
INV_X1 g_I11929 (g6190, I11929);
INV_X1 g_g6649 (I11929, g6649);
INV_X1 g_g6650 (g6213, g6650);
INV_X1 g_I11933 (g5847, I11933);
INV_X1 g_g6651 (I11933, g6651);
INV_X1 g_I11936 (g5918, I11936);
INV_X1 g_g6652 (I11936, g6652);
INV_X1 g_I11939 (g6015, I11939);
INV_X1 g_g6653 (I11939, g6653);
INV_X1 g_I11942 (g6015, I11942);
INV_X1 g_g6654 (I11942, g6654);
INV_X1 g_I11945 (g5874, I11945);
INV_X1 g_g6655 (I11945, g6655);
INV_X1 g_I11948 (g5897, I11948);
INV_X1 g_g6656 (I11948, g6656);
INV_X1 g_I11951 (g5847, I11951);
INV_X1 g_g6657 (I11951, g6657);
INV_X1 g_g6658 (g6224, g6658);
INV_X1 g_I11955 (g5988, I11955);
INV_X1 g_g6659 (I11955, g6659);
INV_X1 g_I11958 (g5874, I11958);
INV_X1 g_g6660 (I11958, g6660);
INV_X1 g_I11961 (g5988, I11961);
INV_X1 g_g6661 (I11961, g6661);
INV_X1 g_I11964 (g5971, I11964);
INV_X1 g_g6662 (I11964, g6662);
INV_X1 g_I11967 (g5971, I11967);
INV_X1 g_g6663 (I11967, g6663);
INV_X1 g_I11971 (g6179, I11971);
INV_X1 g_g6671 (I11971, g6671);
INV_X1 g_I11974 (g5956, I11974);
INV_X1 g_g6672 (I11974, g6672);
INV_X1 g_I11978 (g6186, I11978);
INV_X1 g_g6674 (I11978, g6674);
INV_X1 g_I11981 (g6246, I11981);
INV_X1 g_g6675 (I11981, g6675);
INV_X1 g_I11984 (g6246, I11984);
INV_X1 g_g6676 (I11984, g6676);
INV_X1 g_I11987 (g6278, I11987);
INV_X1 g_g6677 (I11987, g6677);
INV_X1 g_I11991 (g5939, I11991);
INV_X1 g_g6681 (I11991, g6681);
INV_X1 g_I11994 (g6195, I11994);
INV_X1 g_g6682 (I11994, g6682);
INV_X1 g_g6683 (g6237, g6683);
INV_X1 g_I11998 (g5918, I11998);
INV_X1 g_g6684 (I11998, g6684);
INV_X1 g_I12003 (g6202, I12003);
INV_X1 g_g6687 (I12003, g6687);
INV_X1 g_I12008 (g5897, I12008);
INV_X1 g_g6692 (I12008, g6692);
INV_X1 g_I12011 (g5939, I12011);
INV_X1 g_g6693 (I12011, g6693);
INV_X1 g_I12022 (g5874, I12022);
INV_X1 g_g6696 (I12022, g6696);
INV_X1 g_I12025 (g5918, I12025);
INV_X1 g_g6697 (I12025, g6697);
INV_X1 g_g6700 (g6244, g6700);
INV_X1 g_I12038 (g5847, I12038);
INV_X1 g_g6702 (I12038, g6702);
INV_X1 g_I12041 (g5897, I12041);
INV_X1 g_g6703 (I12041, g6703);
INV_X1 g_I12044 (g5847, I12044);
INV_X1 g_g6704 (I12044, g6704);
INV_X1 g_g6708 (g6250, g6708);
INV_X1 g_I12059 (g5874, I12059);
INV_X1 g_g6711 (I12059, g6711);
INV_X1 g_I12062 (g5988, I12062);
INV_X1 g_g6712 (I12062, g6712);
INV_X1 g_I12065 (g5897, I12065);
INV_X1 g_g6713 (I12065, g6713);
INV_X1 g_I12068 (g5847, I12068);
INV_X1 g_g6714 (I12068, g6714);
INV_X1 g_g6720 (g6254, g6720);
INV_X1 g_g6721 (g6257, g6721);
INV_X1 g_I12085 (g5971, I12085);
INV_X1 g_g6723 (I12085, g6723);
INV_X1 g_I12088 (g5874, I12088);
INV_X1 g_g6724 (I12088, g6724);
INV_X1 g_I12091 (g5988, I12091);
INV_X1 g_g6725 (I12091, g6725);
INV_X1 g_g6729 (g6263, g6729);
INV_X1 g_I12098 (g5956, I12098);
INV_X1 g_g6730 (I12098, g6730);
INV_X1 g_I12101 (g5971, I12101);
INV_X1 g_g6731 (I12101, g6731);
INV_X1 g_I12108 (g5939, I12108);
INV_X1 g_g6736 (I12108, g6736);
INV_X1 g_I12111 (g5956, I12111);
INV_X1 g_g6737 (I12111, g6737);
INV_X1 g_I12117 (g5918, I12117);
INV_X1 g_g6741 (I12117, g6741);
INV_X1 g_I12120 (g5939, I12120);
INV_X1 g_g6742 (I12120, g6742);
INV_X1 g_I12124 (g5847, I12124);
INV_X1 g_g6744 (I12124, g6744);
INV_X1 g_I12128 (g5897, I12128);
INV_X1 g_g6751 (I12128, g6751);
INV_X1 g_I12131 (g5918, I12131);
INV_X1 g_g6752 (I12131, g6752);
INV_X1 g_I12135 (g5988, I12135);
INV_X1 g_g6754 (I12135, g6754);
INV_X1 g_I12138 (g5874, I12138);
INV_X1 g_g6755 (I12138, g6755);
INV_X1 g_I12141 (g5897, I12141);
INV_X1 g_g6756 (I12141, g6756);
INV_X1 g_I12145 (g5971, I12145);
INV_X1 g_g6758 (I12145, g6758);
INV_X1 g_I12148 (g5988, I12148);
INV_X1 g_g6759 (I12148, g6759);
INV_X1 g_I12151 (g5847, I12151);
INV_X1 g_g6760 (I12151, g6760);
INV_X1 g_I12154 (g5874, I12154);
INV_X1 g_g6761 (I12154, g6761);
INV_X1 g_I12158 (g5956, I12158);
INV_X1 g_g6763 (I12158, g6763);
INV_X1 g_I12161 (g5971, I12161);
INV_X1 g_g6764 (I12161, g6764);
INV_X1 g_I12164 (g5847, I12164);
INV_X1 g_g6765 (I12164, g6765);
INV_X1 g_I12167 (g5939, I12167);
INV_X1 g_g6766 (I12167, g6766);
INV_X1 g_I12170 (g5956, I12170);
INV_X1 g_g6767 (I12170, g6767);
INV_X1 g_I12173 (g5918, I12173);
INV_X1 g_g6768 (I12173, g6768);
INV_X1 g_I12176 (g5939, I12176);
INV_X1 g_g6769 (I12176, g6769);
INV_X1 g_I12187 (g5897, I12187);
INV_X1 g_g6772 (I12187, g6772);
INV_X1 g_I12190 (g5918, I12190);
INV_X1 g_g6773 (I12190, g6773);
INV_X1 g_I12193 (g6468, I12193);
INV_X1 g_g6774 (I12193, g6774);
INV_X1 g_I12196 (g6471, I12196);
INV_X1 g_g6775 (I12196, g6775);
INV_X1 g_I12199 (g6475, I12199);
INV_X1 g_g6776 (I12199, g6776);
INV_X1 g_I12202 (g6481, I12202);
INV_X1 g_g6777 (I12202, g6777);
INV_X1 g_I12205 (g6488, I12205);
INV_X1 g_g6778 (I12205, g6778);
INV_X1 g_I12208 (g6496, I12208);
INV_X1 g_g6779 (I12208, g6779);
INV_X1 g_I12211 (g6502, I12211);
INV_X1 g_g6780 (I12211, g6780);
INV_X1 g_I12214 (g6507, I12214);
INV_X1 g_g6781 (I12214, g6781);
INV_X1 g_I12217 (g6631, I12217);
INV_X1 g_g6782 (I12217, g6782);
INV_X1 g_I12220 (g6645, I12220);
INV_X1 g_g6783 (I12220, g6783);
INV_X1 g_I12223 (g6655, I12223);
INV_X1 g_g6784 (I12223, g6784);
INV_X1 g_I12226 (g6636, I12226);
INV_X1 g_g6785 (I12226, g6785);
INV_X1 g_I12229 (g6659, I12229);
INV_X1 g_g6786 (I12229, g6786);
INV_X1 g_I12232 (g6662, I12232);
INV_X1 g_g6787 (I12232, g6787);
INV_X1 g_I12235 (g6634, I12235);
INV_X1 g_g6788 (I12235, g6788);
INV_X1 g_I12238 (g6637, I12238);
INV_X1 g_g6789 (I12238, g6789);
INV_X1 g_I12241 (g6640, I12241);
INV_X1 g_g6790 (I12241, g6790);
INV_X1 g_I12244 (g6642, I12244);
INV_X1 g_g6791 (I12244, g6791);
INV_X1 g_I12247 (g6646, I12247);
INV_X1 g_g6792 (I12247, g6792);
INV_X1 g_I12250 (g6651, I12250);
INV_X1 g_g6793 (I12250, g6793);
INV_X1 g_I12253 (g6427, I12253);
INV_X1 g_g6794 (I12253, g6794);
INV_X1 g_I12256 (g6647, I12256);
INV_X1 g_g6795 (I12256, g6795);
INV_X1 g_I12259 (g6652, I12259);
INV_X1 g_g6796 (I12259, g6796);
INV_X1 g_I12262 (g6656, I12262);
INV_X1 g_g6797 (I12262, g6797);
INV_X1 g_I12265 (g6660, I12265);
INV_X1 g_g6798 (I12265, g6798);
INV_X1 g_I12268 (g6661, I12268);
INV_X1 g_g6799 (I12268, g6799);
INV_X1 g_I12271 (g6663, I12271);
INV_X1 g_g6800 (I12271, g6800);
INV_X1 g_I12274 (g6672, I12274);
INV_X1 g_g6801 (I12274, g6801);
INV_X1 g_I12277 (g6681, I12277);
INV_X1 g_g6802 (I12277, g6802);
INV_X1 g_I12280 (g6684, I12280);
INV_X1 g_g6803 (I12280, g6803);
INV_X1 g_I12283 (g6692, I12283);
INV_X1 g_g6804 (I12283, g6804);
INV_X1 g_I12286 (g6696, I12286);
INV_X1 g_g6805 (I12286, g6805);
INV_X1 g_I12289 (g6702, I12289);
INV_X1 g_g6806 (I12289, g6806);
INV_X1 g_I12292 (g6657, I12292);
INV_X1 g_g6807 (I12292, g6807);
INV_X1 g_I12295 (g6693, I12295);
INV_X1 g_g6808 (I12295, g6808);
INV_X1 g_I12298 (g6697, I12298);
INV_X1 g_g6809 (I12298, g6809);
INV_X1 g_I12301 (g6703, I12301);
INV_X1 g_g6810 (I12301, g6810);
INV_X1 g_I12304 (g6711, I12304);
INV_X1 g_g6811 (I12304, g6811);
INV_X1 g_I12307 (g6712, I12307);
INV_X1 g_g6812 (I12307, g6812);
INV_X1 g_I12310 (g6723, I12310);
INV_X1 g_g6813 (I12310, g6813);
INV_X1 g_I12313 (g6730, I12313);
INV_X1 g_g6814 (I12313, g6814);
INV_X1 g_I12316 (g6736, I12316);
INV_X1 g_g6815 (I12316, g6815);
INV_X1 g_I12319 (g6741, I12319);
INV_X1 g_g6816 (I12319, g6816);
INV_X1 g_I12322 (g6751, I12322);
INV_X1 g_g6817 (I12322, g6817);
INV_X1 g_I12325 (g6755, I12325);
INV_X1 g_g6818 (I12325, g6818);
INV_X1 g_I12328 (g6760, I12328);
INV_X1 g_g6819 (I12328, g6819);
INV_X1 g_I12331 (g6704, I12331);
INV_X1 g_g6820 (I12331, g6820);
INV_X1 g_I12334 (g6713, I12334);
INV_X1 g_g6821 (I12334, g6821);
INV_X1 g_I12337 (g6724, I12337);
INV_X1 g_g6822 (I12337, g6822);
INV_X1 g_I12340 (g6725, I12340);
INV_X1 g_g6823 (I12340, g6823);
INV_X1 g_I12343 (g6731, I12343);
INV_X1 g_g6824 (I12343, g6824);
INV_X1 g_I12346 (g6737, I12346);
INV_X1 g_g6825 (I12346, g6825);
INV_X1 g_I12349 (g6742, I12349);
INV_X1 g_g6826 (I12349, g6826);
INV_X1 g_I12352 (g6752, I12352);
INV_X1 g_g6827 (I12352, g6827);
INV_X1 g_I12355 (g6756, I12355);
INV_X1 g_g6828 (I12355, g6828);
INV_X1 g_I12358 (g6761, I12358);
INV_X1 g_g6829 (I12358, g6829);
INV_X1 g_I12361 (g6765, I12361);
INV_X1 g_g6830 (I12361, g6830);
INV_X1 g_I12364 (g6714, I12364);
INV_X1 g_g6831 (I12364, g6831);
INV_X1 g_I12367 (g6754, I12367);
INV_X1 g_g6832 (I12367, g6832);
INV_X1 g_I12370 (g6758, I12370);
INV_X1 g_g6833 (I12370, g6833);
INV_X1 g_I12373 (g6763, I12373);
INV_X1 g_g6834 (I12373, g6834);
INV_X1 g_I12376 (g6766, I12376);
INV_X1 g_g6835 (I12376, g6835);
INV_X1 g_I12379 (g6768, I12379);
INV_X1 g_g6836 (I12379, g6836);
INV_X1 g_I12382 (g6772, I12382);
INV_X1 g_g6837 (I12382, g6837);
INV_X1 g_I12385 (g6397, I12385);
INV_X1 g_g6838 (I12385, g6838);
INV_X1 g_I12388 (g6403, I12388);
INV_X1 g_g6839 (I12388, g6839);
INV_X1 g_I12391 (g6744, I12391);
INV_X1 g_g6840 (I12391, g6840);
INV_X1 g_I12394 (g6759, I12394);
INV_X1 g_g6841 (I12394, g6841);
INV_X1 g_I12397 (g6764, I12397);
INV_X1 g_g6842 (I12397, g6842);
INV_X1 g_I12400 (g6767, I12400);
INV_X1 g_g6843 (I12400, g6843);
INV_X1 g_I12403 (g6769, I12403);
INV_X1 g_g6844 (I12403, g6844);
INV_X1 g_I12406 (g6773, I12406);
INV_X1 g_g6845 (I12406, g6845);
INV_X1 g_I12409 (g6398, I12409);
INV_X1 g_g6846 (I12409, g6846);
INV_X1 g_I12412 (g6404, I12412);
INV_X1 g_g6847 (I12412, g6847);
INV_X1 g_I12415 (g6410, I12415);
INV_X1 g_g6848 (I12415, g6848);
INV_X1 g_I12418 (g6572, I12418);
INV_X1 g_g6849 (I12418, g6849);
INV_X1 g_I12421 (g6486, I12421);
INV_X1 g_g6850 (I12421, g6850);
INV_X1 g_I12424 (g6446, I12424);
INV_X1 g_g6851 (I12424, g6851);
INV_X1 g_I12427 (g6553, I12427);
INV_X1 g_g6852 (I12427, g6852);
INV_X1 g_I12430 (g6432, I12430);
INV_X1 g_g6853 (I12430, g6853);
INV_X1 g_I12433 (g6632, I12433);
INV_X1 g_g6854 (I12433, g6854);
INV_X1 g_I12436 (g6635, I12436);
INV_X1 g_g6855 (I12436, g6855);
INV_X1 g_I12439 (g6566, I12439);
INV_X1 g_g6856 (I12439, g6856);
INV_X1 g_I12442 (g6542, I12442);
INV_X1 g_g6857 (I12442, g6857);
INV_X1 g_I12445 (g6568, I12445);
INV_X1 g_g6858 (I12445, g6858);
INV_X1 g_I12448 (g6569, I12448);
INV_X1 g_g6859 (I12448, g6859);
INV_X1 g_I12451 (g6524, I12451);
INV_X1 g_g6860 (I12451, g6860);
INV_X1 g_I12454 (g6581, I12454);
INV_X1 g_g6861 (I12454, g6861);
INV_X1 g_I12457 (g6671, I12457);
INV_X1 g_g6862 (I12457, g6862);
INV_X1 g_I12460 (g6674, I12460);
INV_X1 g_g6863 (I12460, g6863);
INV_X1 g_I12463 (g6682, I12463);
INV_X1 g_g6864 (I12463, g6864);
INV_X1 g_I12466 (g6687, I12466);
INV_X1 g_g6865 (I12466, g6865);
INV_X1 g_I12469 (g6586, I12469);
INV_X1 g_g6866 (I12469, g6866);
INV_X1 g_I12472 (g6591, I12472);
INV_X1 g_g6867 (I12472, g6867);
INV_X1 g_I12475 (g6596, I12475);
INV_X1 g_g6868 (I12475, g6868);
INV_X1 g_I12478 (g6603, I12478);
INV_X1 g_g6869 (I12478, g6869);
INV_X1 g_I12481 (g6616, I12481);
INV_X1 g_g6870 (I12481, g6870);
INV_X1 g_I12484 (g6621, I12484);
INV_X1 g_g6871 (I12484, g6871);
INV_X1 g_I12487 (g6623, I12487);
INV_X1 g_g6872 (I12487, g6872);
INV_X1 g_I12490 (g6625, I12490);
INV_X1 g_g6873 (I12490, g6873);
INV_X1 g_I12493 (g6587, I12493);
INV_X1 g_g6874 (I12493, g6874);
INV_X1 g_I12496 (g6592, I12496);
INV_X1 g_g6875 (I12496, g6875);
INV_X1 g_I12499 (g6597, I12499);
INV_X1 g_g6876 (I12499, g6876);
INV_X1 g_I12502 (g6604, I12502);
INV_X1 g_g6877 (I12502, g6877);
INV_X1 g_I12505 (g6612, I12505);
INV_X1 g_g6878 (I12505, g6878);
INV_X1 g_I12508 (g6593, I12508);
INV_X1 g_g6879 (I12508, g6879);
INV_X1 g_I12511 (g6598, I12511);
INV_X1 g_g6880 (I12511, g6880);
INV_X1 g_I12514 (g6605, I12514);
INV_X1 g_g6881 (I12514, g6881);
INV_X1 g_I12517 (g6613, I12517);
INV_X1 g_g6882 (I12517, g6882);
INV_X1 g_I12520 (g6622, I12520);
INV_X1 g_g6883 (I12520, g6883);
INV_X1 g_I12523 (g6624, I12523);
INV_X1 g_g6884 (I12523, g6884);
INV_X1 g_I12526 (g6626, I12526);
INV_X1 g_g6885 (I12526, g6885);
INV_X1 g_I12529 (g6628, I12529);
INV_X1 g_g6886 (I12529, g6886);
INV_X1 g_I12532 (g6594, I12532);
INV_X1 g_g6887 (I12532, g6887);
INV_X1 g_I12535 (g6599, I12535);
INV_X1 g_g6888 (I12535, g6888);
INV_X1 g_I12538 (g6606, I12538);
INV_X1 g_g6889 (I12538, g6889);
INV_X1 g_I12541 (g6614, I12541);
INV_X1 g_g6890 (I12541, g6890);
INV_X1 g_I12544 (g6617, I12544);
INV_X1 g_g6891 (I12544, g6891);
INV_X1 g_I12547 (g6708, I12547);
INV_X1 g_g6892 (I12547, g6892);
INV_X1 g_g6894 (g6525, g6894);
INV_X1 g_I12558 (g6449, I12558);
INV_X1 g_g6895 (I12558, g6895);
INV_X1 g_I12561 (g6449, I12561);
INV_X1 g_g6896 (I12561, g6896);
INV_X1 g_I12564 (g6720, I12564);
INV_X1 g_g6897 (I12564, g6897);
INV_X1 g_I12567 (g6721, I12567);
INV_X1 g_g6898 (I12567, g6898);
INV_X1 g_g6899 (g6525, g6899);
INV_X1 g_I12571 (g6729, I12571);
INV_X1 g_g6900 (I12571, g6900);
INV_X1 g_g6901 (g6525, g6901);
INV_X1 g_I12582 (g6745, I12582);
INV_X1 g_g6903 (I12582, g6903);
INV_X1 g_g6904 (g6426, g6904);
INV_X1 g_I12586 (g6643, I12586);
INV_X1 g_g6905 (I12586, g6905);
INV_X1 g_I12592 (g1008, I12592);
INV_X1 g_g6909 (I12592, g6909);
INV_X1 g_I12609 (g6571, I12609);
INV_X1 g_g6918 (I12609, g6918);
INV_X1 g_g6922 (g6525, g6922);
INV_X1 g_I12629 (g6523, I12629);
INV_X1 g_g6936 (I12629, g6936);
INV_X1 g_I12632 (g6514, I12632);
INV_X1 g_g6937 (I12632, g6937);
INV_X1 g_I12635 (g6509, I12635);
INV_X1 g_g6938 (I12635, g6938);
INV_X1 g_g6939 (g6543, g6939);
INV_X1 g_I12639 (g6506, I12639);
INV_X1 g_g6940 (I12639, g6940);
INV_X1 g_I12643 (g6501, I12643);
INV_X1 g_g6944 (I12643, g6944);
INV_X1 g_I12646 (g6493, I12646);
INV_X1 g_g6945 (I12646, g6945);
INV_X1 g_I12649 (g6457, I12649);
INV_X1 g_g6946 (I12649, g6946);
INV_X1 g_I12652 (g6664, I12652);
INV_X1 g_g6947 (I12652, g6947);
INV_X1 g_I12655 (g6458, I12655);
INV_X1 g_g6948 (I12655, g6948);
INV_X1 g_I12659 (g6459, I12659);
INV_X1 g_g6950 (I12659, g6950);
INV_X1 g_g6953 (g6745, g6953);
INV_X1 g_I12666 (g6476, I12666);
INV_X1 g_g6955 (I12666, g6955);
INV_X1 g_I12669 (g6477, I12669);
INV_X1 g_g6956 (I12669, g6956);
INV_X1 g_I12672 (g6473, I12672);
INV_X1 g_g6957 (I12672, g6957);
INV_X1 g_I12675 (g6510, I12675);
INV_X1 g_g6958 (I12675, g6958);
INV_X1 g_I12678 (g6516, I12678);
INV_X1 g_g6959 (I12678, g6959);
INV_X1 g_I12681 (g6469, I12681);
INV_X1 g_g6960 (I12681, g6960);
INV_X1 g_I12684 (g6472, I12684);
INV_X1 g_g6961 (I12684, g6961);
INV_X1 g_I12687 (g6745, I12687);
INV_X1 g_g6962 (I12687, g6962);
INV_X1 g_I12690 (g6467, I12690);
INV_X1 g_g6963 (I12690, g6963);
INV_X1 g_I12696 (g6503, I12696);
INV_X1 g_g6967 (I12696, g6967);
INV_X1 g_I12699 (g6504, I12699);
INV_X1 g_g6968 (I12699, g6968);
INV_X1 g_I12702 (g6497, I12702);
INV_X1 g_g6969 (I12702, g6969);
INV_X1 g_I12708 (g6482, I12708);
INV_X1 g_g6973 (I12708, g6973);
INV_X1 g_I12712 (g6543, I12712);
INV_X1 g_g6975 (I12712, g6975);
INV_X1 g_g6977 (g6664, g6977);
INV_X1 g_I12717 (g6543, I12717);
INV_X1 g_g6978 (I12717, g6978);
INV_X1 g_I12722 (g6611, I12722);
INV_X1 g_g6983 (I12722, g6983);
INV_X1 g_I12725 (g6565, I12725);
INV_X1 g_g6984 (I12725, g6984);
INV_X1 g_I12731 (g6579, I12731);
INV_X1 g_g6993 (I12731, g6993);
INV_X1 g_I12737 (g6460, I12737);
INV_X1 g_g6997 (I12737, g6997);
INV_X1 g_I12742 (g6590, I12742);
INV_X1 g_g7000 (I12742, g7000);
INV_X1 g_I12748 (g6585, I12748);
INV_X1 g_g7006 (I12748, g7006);
INV_X1 g_I12753 (g6445, I12753);
INV_X1 g_g7009 (I12753, g7009);
INV_X1 g_I12757 (g6577, I12757);
INV_X1 g_g7013 (I12757, g7013);
INV_X1 g_I12760 (g6685, I12760);
INV_X1 g_g7014 (I12760, g7014);
INV_X1 g_I12763 (g6686, I12763);
INV_X1 g_g7015 (I12763, g7015);
INV_X1 g_I12768 (g6718, I12768);
INV_X1 g_g7018 (I12768, g7018);
INV_X1 g_I12771 (g6735, I12771);
INV_X1 g_g7019 (I12771, g7019);
INV_X1 g_I12776 (g6739, I12776);
INV_X1 g_g7022 (I12776, g7022);
INV_X1 g_I12779 (g6740, I12779);
INV_X1 g_g7023 (I12779, g7023);
INV_X1 g_I12782 (g6463, I12782);
INV_X1 g_g7024 (I12782, g7024);
INV_X1 g_g7028 (g6525, g7028);
INV_X1 g_g7032 (g6525, g7032);
INV_X1 g_g7034 (g6525, g7034);
INV_X1 g_g7035 (g6543, g7035);
INV_X1 g_g7037 (g6525, g7037);
INV_X1 g_g7039 (g6543, g7039);
INV_X1 g_g7042 (g6543, g7042);
INV_X1 g_g7043 (g6543, g7043);
INV_X1 g_g7044 (g6543, g7044);
INV_X1 g_g7045 (g6490, g7045);
INV_X1 g_I12806 (g6602, I12806);
INV_X1 g_g7046 (I12806, g7046);
INV_X1 g_g7047 (g6498, g7047);
INV_X1 g_I12810 (g6607, I12810);
INV_X1 g_g7048 (I12810, g7048);
INV_X1 g_I12813 (g6607, I12813);
INV_X1 g_g7049 (I12813, g7049);
INV_X1 g_g7050 (g6618, g7050);
INV_X1 g_g7054 (g6511, g7054);
INV_X1 g_g7055 (g6517, g7055);
INV_X1 g_g7056 (g6520, g7056);
INV_X1 g_g7057 (g6644, g7057);
INV_X1 g_g7058 (g6649, g7058);
INV_X1 g_g7059 (g6538, g7059);
INV_X1 g_g7060 (g6654, g7060);
INV_X1 g_g7061 (g6650, g7061);
INV_X1 g_I12826 (g6441, I12826);
INV_X1 g_g7063 (I12826, g7063);
INV_X1 g_I12829 (g6441, I12829);
INV_X1 g_g7064 (I12829, g7064);
INV_X1 g_I12839 (g6630, I12839);
INV_X1 g_g7066 (I12839, g7066);
INV_X1 g_g7067 (g6658, g7067);
INV_X1 g_g7068 (g6556, g7068);
INV_X1 g_g7070 (g6562, g7070);
INV_X1 g_g7077 (g6676, g7077);
INV_X1 g_g7078 (g6683, g7078);
INV_X1 g_g7090 (g6525, g7090);
INV_X1 g_g7091 (g6525, g7091);
INV_X1 g_I12866 (g6483, I12866);
INV_X1 g_g7092 (I12866, g7092);
INV_X1 g_g7094 (g6525, g7094);
INV_X1 g_I12877 (g6700, I12877);
INV_X1 g_g7095 (I12877, g7095);
INV_X1 g_I12881 (g6478, I12881);
INV_X1 g_g7097 (I12881, g7097);
INV_X1 g_g7098 (g6525, g7098);
INV_X1 g_I12885 (g6946, I12885);
INV_X1 g_g7099 (I12885, g7099);
INV_X1 g_I12888 (g6948, I12888);
INV_X1 g_g7100 (I12888, g7100);
INV_X1 g_I12891 (g6950, I12891);
INV_X1 g_g7101 (I12891, g7101);
INV_X1 g_I12894 (g7009, I12894);
INV_X1 g_g7102 (I12894, g7102);
INV_X1 g_I12897 (g6962, I12897);
INV_X1 g_g7103 (I12897, g7103);
INV_X1 g_I12900 (g6947, I12900);
INV_X1 g_g7104 (I12900, g7104);
INV_X1 g_I12903 (g6905, I12903);
INV_X1 g_g7105 (I12903, g7105);
INV_X1 g_I12906 (g6918, I12906);
INV_X1 g_g7106 (I12906, g7106);
INV_X1 g_I12909 (g7046, I12909);
INV_X1 g_g7107 (I12909, g7107);
INV_X1 g_I12912 (g7006, I12912);
INV_X1 g_g7108 (I12912, g7108);
INV_X1 g_I12915 (g7000, I12915);
INV_X1 g_g7109 (I12915, g7109);
INV_X1 g_I12918 (g7013, I12918);
INV_X1 g_g7110 (I12918, g7110);
INV_X1 g_I12921 (g6993, I12921);
INV_X1 g_g7111 (I12921, g7111);
INV_X1 g_I12924 (g6983, I12924);
INV_X1 g_g7112 (I12924, g7112);
INV_X1 g_I12927 (g7014, I12927);
INV_X1 g_g7113 (I12927, g7113);
INV_X1 g_I12930 (g7019, I12930);
INV_X1 g_g7114 (I12930, g7114);
INV_X1 g_I12933 (g7018, I12933);
INV_X1 g_g7115 (I12933, g7115);
INV_X1 g_I12936 (g7015, I12936);
INV_X1 g_g7116 (I12936, g7116);
INV_X1 g_I12939 (g7022, I12939);
INV_X1 g_g7117 (I12939, g7117);
INV_X1 g_I12942 (g7023, I12942);
INV_X1 g_g7118 (I12942, g7118);
INV_X1 g_I12945 (g7066, I12945);
INV_X1 g_g7119 (I12945, g7119);
INV_X1 g_I12948 (g6919, I12948);
INV_X1 g_g7120 (I12948, g7120);
INV_X1 g_I12958 (g6920, I12958);
INV_X1 g_g7122 (I12958, g7122);
INV_X1 g_I12961 (g6921, I12961);
INV_X1 g_g7123 (I12961, g7123);
INV_X1 g_g7124 (g6896, g7124);
INV_X1 g_I12965 (g6924, I12965);
INV_X1 g_g7125 (I12965, g7125);
INV_X1 g_I12968 (g6925, I12968);
INV_X1 g_g7126 (I12968, g7126);
INV_X1 g_g7127 (g6974, g7127);
INV_X1 g_I12973 (g6927, I12973);
INV_X1 g_g7129 (I12973, g7129);
INV_X1 g_I12976 (g6928, I12976);
INV_X1 g_g7130 (I12976, g7130);
INV_X1 g_g7131 (g6976, g7131);
INV_X1 g_I12980 (g6929, I12980);
INV_X1 g_g7132 (I12980, g7132);
INV_X1 g_I12983 (g6930, I12983);
INV_X1 g_g7133 (I12983, g7133);
INV_X1 g_I12986 (g6931, I12986);
INV_X1 g_g7134 (I12986, g7134);
INV_X1 g_I12989 (g6932, I12989);
INV_X1 g_g7135 (I12989, g7135);
INV_X1 g_I12993 (g6933, I12993);
INV_X1 g_g7137 (I12993, g7137);
INV_X1 g_I12996 (g6934, I12996);
INV_X1 g_g7138 (I12996, g7138);
INV_X1 g_I12999 (g7029, I12999);
INV_X1 g_g7139 (I12999, g7139);
INV_X1 g_I13009 (g6935, I13009);
INV_X1 g_g7141 (I13009, g7141);
INV_X1 g_I13012 (g7071, I13012);
INV_X1 g_g7142 (I13012, g7142);
INV_X1 g_g7143 (g6996, g7143);
INV_X1 g_I13023 (g7040, I13023);
INV_X1 g_g7145 (I13023, g7145);
INV_X1 g_g7146 (g6998, g7146);
INV_X1 g_g7147 (g6904, g7147);
INV_X1 g_I13028 (g7087, I13028);
INV_X1 g_g7148 (I13028, g7148);
INV_X1 g_I13031 (g6984, I13031);
INV_X1 g_g7149 (I13031, g7149);
INV_X1 g_g7150 (g6952, g7150);
INV_X1 g_I13035 (g6964, I13035);
INV_X1 g_g7151 (I13035, g7151);
INV_X1 g_I13039 (g6961, I13039);
INV_X1 g_g7155 (I13039, g7155);
INV_X1 g_I13042 (g6963, I13042);
INV_X1 g_g7156 (I13042, g7156);
INV_X1 g_I13045 (g6955, I13045);
INV_X1 g_g7157 (I13045, g7157);
INV_X1 g_I13048 (g6956, I13048);
INV_X1 g_g7158 (I13048, g7158);
INV_X1 g_I13051 (g6967, I13051);
INV_X1 g_g7159 (I13051, g7159);
INV_X1 g_I13054 (g6960, I13054);
INV_X1 g_g7160 (I13054, g7160);
INV_X1 g_I13057 (g6968, I13057);
INV_X1 g_g7161 (I13057, g7161);
INV_X1 g_I13060 (g6959, I13060);
INV_X1 g_g7162 (I13060, g7162);
INV_X1 g_I13063 (g6973, I13063);
INV_X1 g_g7163 (I13063, g7163);
INV_X1 g_I13066 (g6957, I13066);
INV_X1 g_g7164 (I13066, g7164);
INV_X1 g_I13072 (g6969, I13072);
INV_X1 g_g7168 (I13072, g7168);
INV_X1 g_I13075 (g6958, I13075);
INV_X1 g_g7169 (I13075, g7169);
INV_X1 g_g7171 (g7071, g7171);
INV_X1 g_g7172 (g7092, g7172);
INV_X1 g_g7173 (g6980, g7173);
INV_X1 g_g7174 (g7097, g7174);
INV_X1 g_I13084 (g7071, I13084);
INV_X1 g_g7176 (I13084, g7176);
INV_X1 g_I13088 (g7045, I13088);
INV_X1 g_g7178 (I13088, g7178);
INV_X1 g_I13092 (g7047, I13092);
INV_X1 g_g7180 (I13092, g7180);
INV_X1 g_I13099 (g7054, I13099);
INV_X1 g_g7185 (I13099, g7185);
INV_X1 g_I13103 (g7055, I13103);
INV_X1 g_g7187 (I13103, g7187);
INV_X1 g_I13106 (g7056, I13106);
INV_X1 g_g7188 (I13106, g7188);
INV_X1 g_I13109 (g7059, I13109);
INV_X1 g_g7189 (I13109, g7189);
INV_X1 g_I13112 (g7021, I13112);
INV_X1 g_g7190 (I13112, g7190);
INV_X1 g_I13118 (g7068, I13118);
INV_X1 g_g7194 (I13118, g7194);
INV_X1 g_I13122 (g7070, I13122);
INV_X1 g_g7196 (I13122, g7196);
INV_X1 g_I13126 (g6949, I13126);
INV_X1 g_g7198 (I13126, g7198);
INV_X1 g_I13131 (g6951, I13131);
INV_X1 g_g7205 (I13131, g7205);
INV_X1 g_I13134 (g7017, I13134);
INV_X1 g_g7206 (I13134, g7206);
INV_X1 g_I13137 (g7027, I13137);
INV_X1 g_g7207 (I13137, g7207);
INV_X1 g_I13140 (g6954, I13140);
INV_X1 g_g7208 (I13140, g7208);
INV_X1 g_I13144 (g7031, I13144);
INV_X1 g_g7210 (I13144, g7210);
INV_X1 g_I13147 (g7024, I13147);
INV_X1 g_g7211 (I13147, g7211);
INV_X1 g_I13152 (g6966, I13152);
INV_X1 g_g7216 (I13152, g7216);
INV_X1 g_I13157 (g6997, I13157);
INV_X1 g_g7221 (I13157, g7221);
INV_X1 g_I13161 (g7080, I13161);
INV_X1 g_g7223 (I13161, g7223);
INV_X1 g_I13164 (g7086, I13164);
INV_X1 g_g7224 (I13164, g7224);
INV_X1 g_g7225 (g6936, g7225);
INV_X1 g_g7226 (g6937, g7226);
INV_X1 g_g7229 (g6938, g7229);
INV_X1 g_I13173 (g7089, I13173);
INV_X1 g_g7231 (I13173, g7231);
INV_X1 g_g7233 (g6940, g7233);
INV_X1 g_g7236 (g6944, g7236);
INV_X1 g_g7239 (g6945, g7239);
INV_X1 g_I13185 (g7020, I13185);
INV_X1 g_g7241 (I13185, g7241);
INV_X1 g_I13189 (g7002, I13189);
INV_X1 g_g7243 (I13189, g7243);
INV_X1 g_I13193 (g7007, I13193);
INV_X1 g_g7245 (I13193, g7245);
INV_X1 g_I13196 (g7008, I13196);
INV_X1 g_g7246 (I13196, g7246);
INV_X1 g_I13199 (g7025, I13199);
INV_X1 g_g7247 (I13199, g7247);
INV_X1 g_I13203 (g7088, I13203);
INV_X1 g_g7251 (I13203, g7251);
INV_X1 g_g7253 (g7049, g7253);
INV_X1 g_I13209 (g6912, I13209);
INV_X1 g_g7255 (I13209, g7255);
INV_X1 g_g7256 (g7058, g7256);
INV_X1 g_g7259 (g7060, g7259);
INV_X1 g_g7260 (g7064, g7260);
INV_X1 g_I13225 (g7095, I13225);
INV_X1 g_g7261 (I13225, g7261);
INV_X1 g_I13228 (g6892, I13228);
INV_X1 g_g7262 (I13228, g7262);
INV_X1 g_I13231 (g6897, I13231);
INV_X1 g_g7263 (I13231, g7263);
INV_X1 g_I13234 (g6898, I13234);
INV_X1 g_g7264 (I13234, g7264);
INV_X1 g_g7265 (g7077, g7265);
INV_X1 g_I13238 (g6900, I13238);
INV_X1 g_g7266 (I13238, g7266);
INV_X1 g_I13241 (g7030, I13241);
INV_X1 g_g7267 (I13241, g7267);
INV_X1 g_I13244 (g7033, I13244);
INV_X1 g_g7268 (I13244, g7268);
INV_X1 g_I13247 (g6906, I13247);
INV_X1 g_g7269 (I13247, g7269);
INV_X1 g_I13250 (g7036, I13250);
INV_X1 g_g7270 (I13250, g7270);
INV_X1 g_I13255 (g7057, I13255);
INV_X1 g_g7273 (I13255, g7273);
INV_X1 g_I13258 (g6907, I13258);
INV_X1 g_g7274 (I13258, g7274);
INV_X1 g_I13261 (g7041, I13261);
INV_X1 g_g7275 (I13261, g7275);
INV_X1 g_I13264 (g7061, I13264);
INV_X1 g_g7276 (I13264, g7276);
INV_X1 g_I13267 (g6913, I13267);
INV_X1 g_g7277 (I13267, g7277);
INV_X1 g_I13271 (g7067, I13271);
INV_X1 g_g7279 (I13271, g7279);
INV_X1 g_I13274 (g6917, I13274);
INV_X1 g_g7280 (I13274, g7280);
INV_X1 g_I13277 (g7078, I13277);
INV_X1 g_g7281 (I13277, g7281);
INV_X1 g_I13281 (g7155, I13281);
INV_X1 g_g7283 (I13281, g7283);
INV_X1 g_I13284 (g7156, I13284);
INV_X1 g_g7284 (I13284, g7284);
INV_X1 g_I13287 (g7157, I13287);
INV_X1 g_g7285 (I13287, g7285);
INV_X1 g_I13290 (g7158, I13290);
INV_X1 g_g7286 (I13290, g7286);
INV_X1 g_I13293 (g7159, I13293);
INV_X1 g_g7287 (I13293, g7287);
INV_X1 g_I13296 (g7161, I13296);
INV_X1 g_g7288 (I13296, g7288);
INV_X1 g_I13299 (g7163, I13299);
INV_X1 g_g7289 (I13299, g7289);
INV_X1 g_I13302 (g7164, I13302);
INV_X1 g_g7290 (I13302, g7290);
INV_X1 g_I13305 (g7168, I13305);
INV_X1 g_g7291 (I13305, g7291);
INV_X1 g_I13308 (g7169, I13308);
INV_X1 g_g7292 (I13308, g7292);
INV_X1 g_I13311 (g7162, I13311);
INV_X1 g_g7293 (I13311, g7293);
INV_X1 g_I13314 (g7160, I13314);
INV_X1 g_g7294 (I13314, g7294);
INV_X1 g_I13317 (g7211, I13317);
INV_X1 g_g7295 (I13317, g7295);
INV_X1 g_I13320 (g7139, I13320);
INV_X1 g_g7296 (I13320, g7296);
INV_X1 g_I13323 (g7145, I13323);
INV_X1 g_g7297 (I13323, g7297);
INV_X1 g_I13326 (g7176, I13326);
INV_X1 g_g7298 (I13326, g7298);
INV_X1 g_I13329 (g7247, I13329);
INV_X1 g_g7299 (I13329, g7299);
INV_X1 g_I13332 (g7241, I13332);
INV_X1 g_g7300 (I13332, g7300);
INV_X1 g_I13335 (g7206, I13335);
INV_X1 g_g7301 (I13335, g7301);
INV_X1 g_I13338 (g7190, I13338);
INV_X1 g_g7302 (I13338, g7302);
INV_X1 g_I13341 (g7207, I13341);
INV_X1 g_g7303 (I13341, g7303);
INV_X1 g_I13344 (g7210, I13344);
INV_X1 g_g7304 (I13344, g7304);
INV_X1 g_I13347 (g7224, I13347);
INV_X1 g_g7305 (I13347, g7305);
INV_X1 g_I13350 (g7223, I13350);
INV_X1 g_g7306 (I13350, g7306);
INV_X1 g_I13353 (g7231, I13353);
INV_X1 g_g7307 (I13353, g7307);
INV_X1 g_I13356 (g7221, I13356);
INV_X1 g_g7308 (I13356, g7308);
INV_X1 g_I13359 (g7255, I13359);
INV_X1 g_g7309 (I13359, g7309);
INV_X1 g_I13362 (g7265, I13362);
INV_X1 g_g7310 (I13362, g7310);
INV_X1 g_I13365 (g7267, I13365);
INV_X1 g_g7311 (I13365, g7311);
INV_X1 g_I13369 (g7268, I13369);
INV_X1 g_g7313 (I13369, g7313);
INV_X1 g_I13373 (g7270, I13373);
INV_X1 g_g7315 (I13373, g7315);
INV_X1 g_I13383 (g7275, I13383);
INV_X1 g_g7317 (I13383, g7317);
INV_X1 g_g7319 (g7124, g7319);
INV_X1 g_I13388 (g7149, I13388);
INV_X1 g_g7320 (I13388, g7320);
INV_X1 g_I13403 (g7269, I13403);
INV_X1 g_g7327 (I13403, g7327);
INV_X1 g_I13407 (g7271, I13407);
INV_X1 g_g7329 (I13407, g7329);
INV_X1 g_I13410 (g7274, I13410);
INV_X1 g_g7330 (I13410, g7330);
INV_X1 g_I13413 (g7127, I13413);
INV_X1 g_g7331 (I13413, g7331);
INV_X1 g_I13416 (g7165, I13416);
INV_X1 g_g7332 (I13416, g7332);
INV_X1 g_I13419 (g7277, I13419);
INV_X1 g_g7333 (I13419, g7333);
INV_X1 g_I13422 (g7131, I13422);
INV_X1 g_g7334 (I13422, g7334);
INV_X1 g_I13425 (g7166, I13425);
INV_X1 g_g7335 (I13425, g7335);
INV_X1 g_I13428 (g7167, I13428);
INV_X1 g_g7336 (I13428, g7336);
INV_X1 g_I13432 (g7280, I13432);
INV_X1 g_g7338 (I13432, g7338);
INV_X1 g_I13435 (g7170, I13435);
INV_X1 g_g7339 (I13435, g7339);
INV_X1 g_I13438 (g7143, I13438);
INV_X1 g_g7340 (I13438, g7340);
INV_X1 g_I13441 (g7146, I13441);
INV_X1 g_g7341 (I13441, g7341);
INV_X1 g_I13444 (g7282, I13444);
INV_X1 g_g7342 (I13444, g7342);
INV_X1 g_I13447 (g7261, I13447);
INV_X1 g_g7343 (I13447, g7343);
INV_X1 g_g7344 (g7150, g7344);
INV_X1 g_I13451 (g7262, I13451);
INV_X1 g_g7345 (I13451, g7345);
INV_X1 g_I13454 (g7147, I13454);
INV_X1 g_g7346 (I13454, g7346);
INV_X1 g_I13457 (g7120, I13457);
INV_X1 g_g7347 (I13457, g7347);
INV_X1 g_I13460 (g7263, I13460);
INV_X1 g_g7348 (I13460, g7348);
INV_X1 g_I13463 (g7264, I13463);
INV_X1 g_g7349 (I13463, g7349);
INV_X1 g_I13466 (g7122, I13466);
INV_X1 g_g7350 (I13466, g7350);
INV_X1 g_I13469 (g7123, I13469);
INV_X1 g_g7351 (I13469, g7351);
INV_X1 g_I13472 (g7266, I13472);
INV_X1 g_g7352 (I13472, g7352);
INV_X1 g_I13475 (g7125, I13475);
INV_X1 g_g7353 (I13475, g7353);
INV_X1 g_I13478 (g7126, I13478);
INV_X1 g_g7354 (I13478, g7354);
INV_X1 g_I13481 (g7254, I13481);
INV_X1 g_g7355 (I13481, g7355);
INV_X1 g_I13484 (g7128, I13484);
INV_X1 g_g7356 (I13484, g7356);
INV_X1 g_I13487 (g7129, I13487);
INV_X1 g_g7357 (I13487, g7357);
INV_X1 g_I13490 (g7130, I13490);
INV_X1 g_g7358 (I13490, g7358);
INV_X1 g_I13493 (g7132, I13493);
INV_X1 g_g7359 (I13493, g7359);
INV_X1 g_I13496 (g7133, I13496);
INV_X1 g_g7360 (I13496, g7360);
INV_X1 g_I13499 (g7134, I13499);
INV_X1 g_g7361 (I13499, g7361);
INV_X1 g_I13502 (g7135, I13502);
INV_X1 g_g7362 (I13502, g7362);
INV_X1 g_I13506 (g7148, I13506);
INV_X1 g_g7364 (I13506, g7364);
INV_X1 g_I13509 (g7137, I13509);
INV_X1 g_g7365 (I13509, g7365);
INV_X1 g_I13512 (g7138, I13512);
INV_X1 g_g7366 (I13512, g7366);
INV_X1 g_I13515 (g7152, I13515);
INV_X1 g_g7367 (I13515, g7367);
INV_X1 g_I13518 (g7141, I13518);
INV_X1 g_g7405 (I13518, g7405);
INV_X1 g_g7411 (g7202, g7411);
INV_X1 g_I13524 (g7151, I13524);
INV_X1 g_g7413 (I13524, g7413);
INV_X1 g_I13527 (g7217, I13527);
INV_X1 g_g7414 (I13527, g7414);
INV_X1 g_I13533 (g7220, I13533);
INV_X1 g_g7418 (I13533, g7418);
INV_X1 g_I13537 (g7152, I13537);
INV_X1 g_g7420 (I13537, g7420);
INV_X1 g_I13541 (g7209, I13541);
INV_X1 g_g7422 (I13541, g7422);
INV_X1 g_I13544 (g1167, I13544);
INV_X1 g_g7423 (I13544, g7423);
INV_X1 g_I13547 (g1170, I13547);
INV_X1 g_g7424 (I13547, g7424);
INV_X1 g_I13550 (g1173, I13550);
INV_X1 g_g7425 (I13550, g7425);
INV_X1 g_I13559 (g7177, I13559);
INV_X1 g_g7432 (I13559, g7432);
INV_X1 g_I13562 (g7179, I13562);
INV_X1 g_g7433 (I13562, g7433);
INV_X1 g_I13565 (g7181, I13565);
INV_X1 g_g7434 (I13565, g7434);
INV_X1 g_I13570 (g7198, I13570);
INV_X1 g_g7437 (I13570, g7437);
INV_X1 g_I13574 (g7205, I13574);
INV_X1 g_g7439 (I13574, g7439);
INV_X1 g_I13577 (g7186, I13577);
INV_X1 g_g7440 (I13577, g7440);
INV_X1 g_I13580 (g7208, I13580);
INV_X1 g_g7441 (I13580, g7441);
INV_X1 g_I13583 (g7252, I13583);
INV_X1 g_g7442 (I13583, g7442);
INV_X1 g_I13595 (g7216, I13595);
INV_X1 g_g7446 (I13595, g7446);
INV_X1 g_I13605 (g7197, I13605);
INV_X1 g_g7448 (I13605, g7448);
INV_X1 g_I13610 (g7227, I13610);
INV_X1 g_g7454 (I13610, g7454);
INV_X1 g_I13613 (g7273, I13613);
INV_X1 g_g7455 (I13613, g7455);
INV_X1 g_g7456 (g7174, g7456);
INV_X1 g_I13617 (g7276, I13617);
INV_X1 g_g7459 (I13617, g7459);
INV_X1 g_g7460 (g7172, g7460);
INV_X1 g_g7463 (g7239, g7463);
INV_X1 g_I13622 (g7279, I13622);
INV_X1 g_g7466 (I13622, g7466);
INV_X1 g_g7467 (g7236, g7467);
INV_X1 g_g7470 (g7253, g7470);
INV_X1 g_g7471 (g7233, g7471);
INV_X1 g_I13628 (g7248, I13628);
INV_X1 g_g7474 (I13628, g7474);
INV_X1 g_I13631 (g7248, I13631);
INV_X1 g_g7475 (I13631, g7475);
INV_X1 g_g7476 (g7229, g7476);
INV_X1 g_I13635 (g7243, I13635);
INV_X1 g_g7479 (I13635, g7479);
INV_X1 g_g7483 (g7226, g7483);
INV_X1 g_I13646 (g7245, I13646);
INV_X1 g_g7486 (I13646, g7486);
INV_X1 g_I13649 (g7281, I13649);
INV_X1 g_g7487 (I13649, g7487);
INV_X1 g_g7488 (g7225, g7488);
INV_X1 g_I13653 (g7246, I13653);
INV_X1 g_g7491 (I13653, g7491);
INV_X1 g_I13656 (g7228, I13656);
INV_X1 g_g7492 (I13656, g7492);
INV_X1 g_I13659 (g7232, I13659);
INV_X1 g_g7493 (I13659, g7493);
INV_X1 g_g7494 (g7260, g7494);
INV_X1 g_I13663 (g7235, I13663);
INV_X1 g_g7495 (I13663, g7495);
INV_X1 g_I13666 (g7238, I13666);
INV_X1 g_g7496 (I13666, g7496);
INV_X1 g_I13669 (g7240, I13669);
INV_X1 g_g7497 (I13669, g7497);
INV_X1 g_I13672 (g7242, I13672);
INV_X1 g_g7498 (I13672, g7498);
INV_X1 g_g7499 (g7258, g7499);
INV_X1 g_I13676 (g7256, I13676);
INV_X1 g_g7500 (I13676, g7500);
INV_X1 g_I13679 (g7259, I13679);
INV_X1 g_g7501 (I13679, g7501);
INV_X1 g_I13682 (g7251, I13682);
INV_X1 g_g7502 (I13682, g7502);
INV_X1 g_I13692 (g7343, I13692);
INV_X1 g_g7504 (I13692, g7504);
INV_X1 g_I13695 (g7345, I13695);
INV_X1 g_g7505 (I13695, g7505);
INV_X1 g_I13698 (g7348, I13698);
INV_X1 g_g7506 (I13698, g7506);
INV_X1 g_I13701 (g7349, I13701);
INV_X1 g_g7507 (I13701, g7507);
INV_X1 g_I13704 (g7352, I13704);
INV_X1 g_g7508 (I13704, g7508);
INV_X1 g_I13707 (g7420, I13707);
INV_X1 g_g7509 (I13707, g7509);
INV_X1 g_I13710 (g7340, I13710);
INV_X1 g_g7510 (I13710, g7510);
INV_X1 g_I13713 (g7341, I13713);
INV_X1 g_g7511 (I13713, g7511);
INV_X1 g_I13716 (g7331, I13716);
INV_X1 g_g7512 (I13716, g7512);
INV_X1 g_I13719 (g7334, I13719);
INV_X1 g_g7513 (I13719, g7513);
INV_X1 g_I13722 (g7442, I13722);
INV_X1 g_g7514 (I13722, g7514);
INV_X1 g_I13725 (g7437, I13725);
INV_X1 g_g7515 (I13725, g7515);
INV_X1 g_I13728 (g7439, I13728);
INV_X1 g_g7516 (I13728, g7516);
INV_X1 g_I13731 (g7441, I13731);
INV_X1 g_g7517 (I13731, g7517);
INV_X1 g_I13734 (g7422, I13734);
INV_X1 g_g7518 (I13734, g7518);
INV_X1 g_I13737 (g7446, I13737);
INV_X1 g_g7519 (I13737, g7519);
INV_X1 g_I13740 (g7364, I13740);
INV_X1 g_g7520 (I13740, g7520);
INV_X1 g_I13743 (g7454, I13743);
INV_X1 g_g7521 (I13743, g7521);
INV_X1 g_I13746 (g7311, I13746);
INV_X1 g_g7522 (I13746, g7522);
INV_X1 g_I13749 (g7313, I13749);
INV_X1 g_g7523 (I13749, g7523);
INV_X1 g_I13752 (g7315, I13752);
INV_X1 g_g7524 (I13752, g7524);
INV_X1 g_I13755 (g7317, I13755);
INV_X1 g_g7525 (I13755, g7525);
INV_X1 g_I13758 (g7414, I13758);
INV_X1 g_g7526 (I13758, g7526);
INV_X1 g_I13761 (g7418, I13761);
INV_X1 g_g7527 (I13761, g7527);
INV_X1 g_I13764 (g7479, I13764);
INV_X1 g_g7528 (I13764, g7528);
INV_X1 g_I13767 (g7486, I13767);
INV_X1 g_g7529 (I13767, g7529);
INV_X1 g_I13770 (g7491, I13770);
INV_X1 g_g7530 (I13770, g7530);
INV_X1 g_I13773 (g7496, I13773);
INV_X1 g_g7531 (I13773, g7531);
INV_X1 g_I13776 (g7497, I13776);
INV_X1 g_g7532 (I13776, g7532);
INV_X1 g_I13779 (g7406, I13779);
INV_X1 g_g7533 (I13779, g7533);
INV_X1 g_I13782 (g7498, I13782);
INV_X1 g_g7534 (I13782, g7534);
INV_X1 g_I13794 (g7346, I13794);
INV_X1 g_g7538 (I13794, g7538);
INV_X1 g_I13797 (g7502, I13797);
INV_X1 g_g7539 (I13797, g7539);
INV_X1 g_I13807 (g7320, I13807);
INV_X1 g_g7541 (I13807, g7541);
INV_X1 g_I13810 (g7312, I13810);
INV_X1 g_g7542 (I13810, g7542);
INV_X1 g_I13813 (g7314, I13813);
INV_X1 g_g7543 (I13813, g7543);
INV_X1 g_I13816 (g7455, I13816);
INV_X1 g_g7544 (I13816, g7544);
INV_X1 g_I13819 (g7426, I13819);
INV_X1 g_g7545 (I13819, g7545);
INV_X1 g_I13822 (g7459, I13822);
INV_X1 g_g7546 (I13822, g7546);
INV_X1 g_I13825 (g7318, I13825);
INV_X1 g_g7547 (I13825, g7547);
INV_X1 g_I13828 (g7321, I13828);
INV_X1 g_g7548 (I13828, g7548);
INV_X1 g_I13831 (g7322, I13831);
INV_X1 g_g7549 (I13831, g7549);
INV_X1 g_I13834 (g7466, I13834);
INV_X1 g_g7550 (I13834, g7550);
INV_X1 g_I13837 (g7324, I13837);
INV_X1 g_g7551 (I13837, g7551);
INV_X1 g_I13843 (g7326, I13843);
INV_X1 g_g7555 (I13843, g7555);
INV_X1 g_I13846 (g7487, I13846);
INV_X1 g_g7556 (I13846, g7556);
INV_X1 g_I13850 (g7328, I13850);
INV_X1 g_g7558 (I13850, g7558);
INV_X1 g_I13854 (g7327, I13854);
INV_X1 g_g7560 (I13854, g7560);
INV_X1 g_I13858 (g7329, I13858);
INV_X1 g_g7562 (I13858, g7562);
INV_X1 g_I13861 (g7330, I13861);
INV_X1 g_g7563 (I13861, g7563);
INV_X1 g_I13865 (g7333, I13865);
INV_X1 g_g7565 (I13865, g7565);
INV_X1 g_I13869 (g7338, I13869);
INV_X1 g_g7574 (I13869, g7574);
INV_X1 g_I13873 (g7342, I13873);
INV_X1 g_g7576 (I13873, g7576);
INV_X1 g_I13876 (g7347, I13876);
INV_X1 g_g7577 (I13876, g7577);
INV_X1 g_I13879 (g7332, I13879);
INV_X1 g_g7578 (I13879, g7578);
INV_X1 g_I13882 (g7350, I13882);
INV_X1 g_g7579 (I13882, g7579);
INV_X1 g_I13885 (g7351, I13885);
INV_X1 g_g7580 (I13885, g7580);
INV_X1 g_I13888 (g7335, I13888);
INV_X1 g_g7581 (I13888, g7581);
INV_X1 g_I13891 (g7336, I13891);
INV_X1 g_g7582 (I13891, g7582);
INV_X1 g_I13894 (g7353, I13894);
INV_X1 g_g7583 (I13894, g7583);
INV_X1 g_I13897 (g7354, I13897);
INV_X1 g_g7584 (I13897, g7584);
INV_X1 g_I13900 (g7356, I13900);
INV_X1 g_g7585 (I13900, g7585);
INV_X1 g_I13903 (g7357, I13903);
INV_X1 g_g7586 (I13903, g7586);
INV_X1 g_I13906 (g7358, I13906);
INV_X1 g_g7587 (I13906, g7587);
INV_X1 g_I13909 (g7339, I13909);
INV_X1 g_g7588 (I13909, g7588);
INV_X1 g_I13912 (g7359, I13912);
INV_X1 g_g7589 (I13912, g7589);
INV_X1 g_I13915 (g7360, I13915);
INV_X1 g_g7590 (I13915, g7590);
INV_X1 g_I13918 (g7361, I13918);
INV_X1 g_g7591 (I13918, g7591);
INV_X1 g_I13921 (g7362, I13921);
INV_X1 g_g7592 (I13921, g7592);
INV_X1 g_I13924 (g7365, I13924);
INV_X1 g_g7593 (I13924, g7593);
INV_X1 g_I13927 (g7366, I13927);
INV_X1 g_g7594 (I13927, g7594);
INV_X1 g_I13930 (g7405, I13930);
INV_X1 g_g7595 (I13930, g7595);
INV_X1 g_g7599 (g7450, g7599);
INV_X1 g_g7601 (g7450, g7601);
INV_X1 g_I13940 (g7355, I13940);
INV_X1 g_g7603 (I13940, g7603);
INV_X1 g_g7610 (g7450, g7610);
INV_X1 g_I13956 (g7499, I13956);
INV_X1 g_g7627 (I13956, g7627);
INV_X1 g_I13962 (g7413, I13962);
INV_X1 g_g7633 (I13962, g7633);
INV_X1 g_I13979 (g7415, I13979);
INV_X1 g_g7686 (I13979, g7686);
INV_X1 g_g7688 (g7406, g7688);
INV_X1 g_I13997 (g7432, I13997);
INV_X1 g_g7702 (I13997, g7702);
INV_X1 g_I14001 (g7433, I14001);
INV_X1 g_g7704 (I14001, g7704);
INV_X1 g_I14005 (g7434, I14005);
INV_X1 g_g7708 (I14005, g7708);
INV_X1 g_I14009 (g7436, I14009);
INV_X1 g_g7710 (I14009, g7710);
INV_X1 g_I14012 (g7438, I14012);
INV_X1 g_g7711 (I14012, g7711);
INV_X1 g_I14015 (g7440, I14015);
INV_X1 g_g7712 (I14015, g7712);
INV_X1 g_I14019 (g7480, I14019);
INV_X1 g_g7714 (I14019, g7714);
INV_X1 g_I14022 (g7443, I14022);
INV_X1 g_g7715 (I14022, g7715);
INV_X1 g_I14025 (g7500, I14025);
INV_X1 g_g7716 (I14025, g7716);
INV_X1 g_I14028 (g7501, I14028);
INV_X1 g_g7717 (I14028, g7717);
INV_X1 g_I14031 (g7448, I14031);
INV_X1 g_g7718 (I14031, g7718);
INV_X1 g_g7719 (g7475, g7719);
INV_X1 g_I14035 (g7310, I14035);
INV_X1 g_g7720 (I14035, g7720);
INV_X1 g_g7721 (g7344, g7721);
INV_X1 g_I14039 (g7449, I14039);
INV_X1 g_g7722 (I14039, g7722);
INV_X1 g_I14042 (g7470, I14042);
INV_X1 g_g7723 (I14042, g7723);
INV_X1 g_I14046 (g7492, I14046);
INV_X1 g_g7725 (I14046, g7725);
INV_X1 g_I14049 (g7493, I14049);
INV_X1 g_g7726 (I14049, g7726);
INV_X1 g_I14052 (g7494, I14052);
INV_X1 g_g7727 (I14052, g7727);
INV_X1 g_I14055 (g7495, I14055);
INV_X1 g_g7728 (I14055, g7728);
INV_X1 g_I14058 (g7544, I14058);
INV_X1 g_g7729 (I14058, g7729);
INV_X1 g_I14061 (g7546, I14061);
INV_X1 g_g7730 (I14061, g7730);
INV_X1 g_I14064 (g7556, I14064);
INV_X1 g_g7731 (I14064, g7731);
INV_X1 g_I14067 (g7550, I14067);
INV_X1 g_g7732 (I14067, g7732);
INV_X1 g_I14070 (g7714, I14070);
INV_X1 g_g7733 (I14070, g7733);
INV_X1 g_I14073 (g7627, I14073);
INV_X1 g_g7734 (I14073, g7734);
INV_X1 g_I14076 (g7577, I14076);
INV_X1 g_g7735 (I14076, g7735);
INV_X1 g_I14079 (g7579, I14079);
INV_X1 g_g7736 (I14079, g7736);
INV_X1 g_I14082 (g7539, I14082);
INV_X1 g_g7737 (I14082, g7737);
INV_X1 g_I14085 (g7583, I14085);
INV_X1 g_g7738 (I14085, g7738);
INV_X1 g_I14088 (g7585, I14088);
INV_X1 g_g7739 (I14088, g7739);
INV_X1 g_I14091 (g7589, I14091);
INV_X1 g_g7740 (I14091, g7740);
INV_X1 g_I14094 (g7593, I14094);
INV_X1 g_g7741 (I14094, g7741);
INV_X1 g_I14097 (g7595, I14097);
INV_X1 g_g7742 (I14097, g7742);
INV_X1 g_I14100 (g7580, I14100);
INV_X1 g_g7743 (I14100, g7743);
INV_X1 g_I14103 (g7584, I14103);
INV_X1 g_g7744 (I14103, g7744);
INV_X1 g_I14106 (g7586, I14106);
INV_X1 g_g7745 (I14106, g7745);
INV_X1 g_I14109 (g7590, I14109);
INV_X1 g_g7746 (I14109, g7746);
INV_X1 g_I14112 (g7560, I14112);
INV_X1 g_g7747 (I14112, g7747);
INV_X1 g_I14115 (g7563, I14115);
INV_X1 g_g7748 (I14115, g7748);
INV_X1 g_I14118 (g7565, I14118);
INV_X1 g_g7749 (I14118, g7749);
INV_X1 g_I14121 (g7587, I14121);
INV_X1 g_g7750 (I14121, g7750);
INV_X1 g_I14124 (g7591, I14124);
INV_X1 g_g7751 (I14124, g7751);
INV_X1 g_I14127 (g7594, I14127);
INV_X1 g_g7752 (I14127, g7752);
INV_X1 g_I14130 (g7592, I14130);
INV_X1 g_g7753 (I14130, g7753);
INV_X1 g_I14133 (g7574, I14133);
INV_X1 g_g7754 (I14133, g7754);
INV_X1 g_I14136 (g7633, I14136);
INV_X1 g_g7755 (I14136, g7755);
INV_X1 g_I14139 (g7548, I14139);
INV_X1 g_g7756 (I14139, g7756);
INV_X1 g_I14142 (g7551, I14142);
INV_X1 g_g7757 (I14142, g7757);
INV_X1 g_I14145 (g7542, I14145);
INV_X1 g_g7758 (I14145, g7758);
INV_X1 g_I14148 (g7543, I14148);
INV_X1 g_g7759 (I14148, g7759);
INV_X1 g_I14151 (g7555, I14151);
INV_X1 g_g7760 (I14151, g7760);
INV_X1 g_I14154 (g7558, I14154);
INV_X1 g_g7761 (I14154, g7761);
INV_X1 g_I14157 (g7547, I14157);
INV_X1 g_g7762 (I14157, g7762);
INV_X1 g_I14160 (g7549, I14160);
INV_X1 g_g7763 (I14160, g7763);
INV_X1 g_I14163 (g7533, I14163);
INV_X1 g_g7764 (I14163, g7764);
INV_X1 g_I14166 (g7702, I14166);
INV_X1 g_g7765 (I14166, g7765);
INV_X1 g_I14169 (g7715, I14169);
INV_X1 g_g7766 (I14169, g7766);
INV_X1 g_I14172 (g7545, I14172);
INV_X1 g_g7767 (I14172, g7767);
INV_X1 g_I14175 (g7718, I14175);
INV_X1 g_g7768 (I14175, g7768);
INV_X1 g_I14178 (g7562, I14178);
INV_X1 g_g7769 (I14178, g7769);
INV_X1 g_I14181 (g7725, I14181);
INV_X1 g_g7770 (I14181, g7770);
INV_X1 g_I14184 (g7726, I14184);
INV_X1 g_g7771 (I14184, g7771);
INV_X1 g_I14187 (g7728, I14187);
INV_X1 g_g7772 (I14187, g7772);
INV_X1 g_I14190 (g7531, I14190);
INV_X1 g_g7773 (I14190, g7773);
INV_X1 g_I14193 (g7532, I14193);
INV_X1 g_g7774 (I14193, g7774);
INV_X1 g_I14196 (g7534, I14196);
INV_X1 g_g7775 (I14196, g7775);
INV_X1 g_I14199 (g7704, I14199);
INV_X1 g_g7776 (I14199, g7776);
INV_X1 g_I14202 (g7708, I14202);
INV_X1 g_g7777 (I14202, g7777);
INV_X1 g_I14205 (g7710, I14205);
INV_X1 g_g7778 (I14205, g7778);
INV_X1 g_I14208 (g7711, I14208);
INV_X1 g_g7779 (I14208, g7779);
INV_X1 g_I14211 (g7712, I14211);
INV_X1 g_g7780 (I14211, g7780);
INV_X1 g_I14214 (g7576, I14214);
INV_X1 g_g7781 (I14214, g7781);
INV_X1 g_I14224 (g7722, I14224);
INV_X1 g_g7789 (I14224, g7789);
INV_X1 g_I14227 (g7552, I14227);
INV_X1 g_g7790 (I14227, g7790);
INV_X1 g_I14231 (g7566, I14231);
INV_X1 g_g7792 (I14231, g7792);
INV_X1 g_I14234 (g7614, I14234);
INV_X1 g_g7793 (I14234, g7793);
INV_X1 g_I14238 (g7608, I14238);
INV_X1 g_g7811 (I14238, g7811);
INV_X1 g_I14251 (g7541, I14251);
INV_X1 g_g7829 (I14251, g7829);
INV_X1 g_I14257 (g7716, I14257);
INV_X1 g_g7835 (I14257, g7835);
INV_X1 g_I14260 (g7717, I14260);
INV_X1 g_g7836 (I14260, g7836);
INV_X1 g_I14264 (g7698, I14264);
INV_X1 g_g7838 (I14264, g7838);
INV_X1 g_I14267 (g7695, I14267);
INV_X1 g_g7855 (I14267, g7855);
INV_X1 g_I14270 (g7703, I14270);
INV_X1 g_g7870 (I14270, g7870);
INV_X1 g_I14273 (g7631, I14273);
INV_X1 g_g7887 (I14273, g7887);
INV_X1 g_I14276 (g7720, I14276);
INV_X1 g_g7904 (I14276, g7904);
INV_X1 g_I14279 (g7700, I14279);
INV_X1 g_g7905 (I14279, g7905);
INV_X1 g_I14282 (g7709, I14282);
INV_X1 g_g7920 (I14282, g7920);
INV_X1 g_I14285 (g7625, I14285);
INV_X1 g_g7937 (I14285, g7937);
INV_X1 g_I14288 (g7705, I14288);
INV_X1 g_g7951 (I14288, g7951);
INV_X1 g_I14291 (g7680, I14291);
INV_X1 g_g7966 (I14291, g7966);
INV_X1 g_I14294 (g7553, I14294);
INV_X1 g_g7983 (I14294, g7983);
INV_X1 g_g7992 (g7557, g7992);
INV_X1 g_I14298 (g7678, I14298);
INV_X1 g_g7993 (I14298, g7993);
INV_X1 g_g8008 (g7559, g8008);
INV_X1 g_I14305 (g7537, I14305);
INV_X1 g_g8012 (I14305, g8012);
INV_X1 g_g8013 (g7561, g8013);
INV_X1 g_g8014 (g7564, g8014);
INV_X1 g_g8015 (g7689, g8015);
INV_X1 g_I14311 (g7566, I14311);
INV_X1 g_g8016 (I14311, g8016);
INV_X1 g_g8017 (g7692, g8017);
INV_X1 g_I14315 (g7676, I14315);
INV_X1 g_g8018 (I14315, g8018);
INV_X1 g_I14318 (g7657, I14318);
INV_X1 g_g8029 (I14318, g8029);
INV_X1 g_g8038 (g7694, g8038);
INV_X1 g_g8039 (g7696, g8039);
INV_X1 g_g8040 (g7699, g8040);
INV_X1 g_g8041 (g7701, g8041);
INV_X1 g_I14325 (g7713, I14325);
INV_X1 g_g8042 (I14325, g8042);
INV_X1 g_I14330 (g7538, I14330);
INV_X1 g_g8061 (I14330, g8061);
INV_X1 g_I14334 (g7578, I14334);
INV_X1 g_g8063 (I14334, g8063);
INV_X1 g_I14338 (g7581, I14338);
INV_X1 g_g8065 (I14338, g8065);
INV_X1 g_I14342 (g7582, I14342);
INV_X1 g_g8067 (I14342, g8067);
INV_X1 g_I14349 (g7588, I14349);
INV_X1 g_g8072 (I14349, g8072);
INV_X1 g_I14370 (g7603, I14370);
INV_X1 g_g8093 (I14370, g8093);
INV_X1 g_g8094 (g7705, g8094);
INV_X1 g_I14374 (g7693, I14374);
INV_X1 g_g8111 (I14374, g8111);
INV_X1 g_I14378 (g7691, I14378);
INV_X1 g_g8131 (I14378, g8131);
INV_X1 g_I14381 (g7596, I14381);
INV_X1 g_g8145 (I14381, g8145);
INV_X1 g_I14388 (g7605, I14388);
INV_X1 g_g8152 (I14388, g8152);
INV_X1 g_I14394 (g7536, I14394);
INV_X1 g_g8156 (I14394, g8156);
INV_X1 g_I14397 (g7686, I14397);
INV_X1 g_g8172 (I14397, g8172);
INV_X1 g_I14400 (g7677, I14400);
INV_X1 g_g8173 (I14400, g8173);
INV_X1 g_I14403 (g7679, I14403);
INV_X1 g_g8174 (I14403, g8174);
INV_X1 g_I14406 (g7681, I14406);
INV_X1 g_g8175 (I14406, g8175);
INV_X1 g_I14410 (g7697, I14410);
INV_X1 g_g8177 (I14410, g8177);
INV_X1 g_I14413 (g7723, I14413);
INV_X1 g_g8178 (I14413, g8178);
INV_X1 g_I14416 (g7727, I14416);
INV_X1 g_g8179 (I14416, g8179);
INV_X1 g_g8180 (g7719, g8180);
INV_X1 g_I14420 (g7554, I14420);
INV_X1 g_g8181 (I14420, g8181);
INV_X1 g_g8198 (g7721, g8198);
INV_X1 g_I14424 (g7652, I14424);
INV_X1 g_g8199 (I14424, g8199);
INV_X1 g_I14427 (g7835, I14427);
INV_X1 g_g8216 (I14427, g8216);
INV_X1 g_I14430 (g7836, I14430);
INV_X1 g_g8217 (I14430, g8217);
INV_X1 g_I14433 (g8061, I14433);
INV_X1 g_g8218 (I14433, g8218);
INV_X1 g_I14436 (g7904, I14436);
INV_X1 g_g8219 (I14436, g8219);
INV_X1 g_I14439 (g8063, I14439);
INV_X1 g_g8220 (I14439, g8220);
INV_X1 g_I14442 (g8065, I14442);
INV_X1 g_g8221 (I14442, g8221);
INV_X1 g_I14445 (g8067, I14445);
INV_X1 g_g8222 (I14445, g8222);
INV_X1 g_I14448 (g7792, I14448);
INV_X1 g_g8223 (I14448, g8223);
INV_X1 g_I14451 (g8172, I14451);
INV_X1 g_g8224 (I14451, g8224);
INV_X1 g_I14454 (g8177, I14454);
INV_X1 g_g8225 (I14454, g8225);
INV_X1 g_I14457 (g8093, I14457);
INV_X1 g_g8226 (I14457, g8226);
INV_X1 g_I14460 (g7789, I14460);
INV_X1 g_g8227 (I14460, g8227);
INV_X1 g_I14463 (g8072, I14463);
INV_X1 g_g8228 (I14463, g8228);
INV_X1 g_I14489 (g7829, I14489);
INV_X1 g_g8234 (I14489, g8234);
INV_X1 g_I14492 (g7829, I14492);
INV_X1 g_g8235 (I14492, g8235);
INV_X1 g_I14531 (g8178, I14531);
INV_X1 g_g8284 (I14531, g8284);
INV_X1 g_I14573 (g8179, I14573);
INV_X1 g_g8324 (I14573, g8324);
INV_X1 g_g8342 (g8008, g8342);
INV_X1 g_g8363 (g7992, g8363);
INV_X1 g_I14603 (g7827, I14603);
INV_X1 g_g8381 (I14603, g8381);
INV_X1 g_g8386 (g8014, g8386);
INV_X1 g_I14614 (g7832, I14614);
INV_X1 g_g8406 (I14614, g8406);
INV_X1 g_g8407 (g8013, g8407);
INV_X1 g_g8421 (g8017, g8421);
INV_X1 g_I14623 (g7833, I14623);
INV_X1 g_g8442 (I14623, g8442);
INV_X1 g_g8443 (g8015, g8443);
INV_X1 g_g8463 (g8094, g8463);
INV_X1 g_g8464 (g8039, g8464);
INV_X1 g_I14637 (g8012, I14637);
INV_X1 g_g8481 (I14637, g8481);
INV_X1 g_g8482 (g8094, g8482);
INV_X1 g_g8483 (g8038, g8483);
INV_X1 g_g8493 (g8041, g8493);
INV_X1 g_I14643 (g7837, I14643);
INV_X1 g_g8510 (I14643, g8510);
INV_X1 g_I14646 (g7790, I14646);
INV_X1 g_g8511 (I14646, g8511);
INV_X1 g_g8512 (g8094, g8512);
INV_X1 g_g8514 (g8040, g8514);
INV_X1 g_g8524 (g7855, g8524);
INV_X1 g_g8541 (g8094, g8541);
INV_X1 g_I14657 (g7782, I14657);
INV_X1 g_g8544 (I14657, g8544);
INV_X1 g_g8545 (g7905, g8545);
INV_X1 g_g8562 (g8094, g8562);
INV_X1 g_I14662 (g7783, I14662);
INV_X1 g_g8563 (I14662, g8563);
INV_X1 g_g8564 (g7951, g8564);
INV_X1 g_g8581 (g8094, g8581);
INV_X1 g_g8582 (g8094, g8582);
INV_X1 g_I14668 (g7787, I14668);
INV_X1 g_g8583 (I14668, g8583);
INV_X1 g_g8585 (g7993, g8585);
INV_X1 g_g8602 (g8094, g8602);
INV_X1 g_I14674 (g7788, I14674);
INV_X1 g_g8603 (I14674, g8603);
INV_X1 g_I14677 (g7791, I14677);
INV_X1 g_g8604 (I14677, g8604);
INV_X1 g_I14680 (g7810, I14680);
INV_X1 g_g8605 (I14680, g8605);
INV_X1 g_I14683 (g7825, I14683);
INV_X1 g_g8606 (I14683, g8606);
INV_X1 g_I14687 (g7826, I14687);
INV_X1 g_g8608 (I14687, g8608);
INV_X1 g_I14695 (g8016, I14695);
INV_X1 g_g8619 (I14695, g8619);
INV_X1 g_I14709 (g8198, I14709);
INV_X1 g_g8631 (I14709, g8631);
INV_X1 g_I14712 (g8059, I14712);
INV_X1 g_g8632 (I14712, g8632);
INV_X1 g_I14718 (g8068, I14718);
INV_X1 g_g8636 (I14718, g8636);
INV_X1 g_I14722 (g8076, I14722);
INV_X1 g_g8638 (I14722, g8638);
INV_X1 g_I14725 (g8145, I14725);
INV_X1 g_g8639 (I14725, g8639);
INV_X1 g_I14728 (g8152, I14728);
INV_X1 g_g8640 (I14728, g8640);
INV_X1 g_I14732 (g8155, I14732);
INV_X1 g_g8642 (I14732, g8642);
INV_X1 g_I14739 (g8173, I14739);
INV_X1 g_g8647 (I14739, g8647);
INV_X1 g_I14743 (g8174, I14743);
INV_X1 g_g8649 (I14743, g8649);
INV_X1 g_I14747 (g8175, I14747);
INV_X1 g_g8651 (I14747, g8651);
INV_X1 g_I14763 (g7834, I14763);
INV_X1 g_g8657 (I14763, g8657);
INV_X1 g_I14777 (g8511, I14777);
INV_X1 g_g8661 (I14777, g8661);
INV_X1 g_I14780 (g8284, I14780);
INV_X1 g_g8662 (I14780, g8662);
INV_X1 g_I14783 (g8324, I14783);
INV_X1 g_g8663 (I14783, g8663);
INV_X1 g_I14786 (g8606, I14786);
INV_X1 g_g8664 (I14786, g8664);
INV_X1 g_I14789 (g8544, I14789);
INV_X1 g_g8665 (I14789, g8665);
INV_X1 g_I14792 (g8583, I14792);
INV_X1 g_g8666 (I14792, g8666);
INV_X1 g_I14795 (g8604, I14795);
INV_X1 g_g8667 (I14795, g8667);
INV_X1 g_I14798 (g8605, I14798);
INV_X1 g_g8668 (I14798, g8668);
INV_X1 g_I14801 (g8608, I14801);
INV_X1 g_g8669 (I14801, g8669);
INV_X1 g_I14804 (g8563, I14804);
INV_X1 g_g8670 (I14804, g8670);
INV_X1 g_I14807 (g8603, I14807);
INV_X1 g_g8671 (I14807, g8671);
INV_X1 g_I14810 (g8481, I14810);
INV_X1 g_g8672 (I14810, g8672);
INV_X1 g_I14813 (g8640, I14813);
INV_X1 g_g8673 (I14813, g8673);
INV_X1 g_I14816 (g8642, I14816);
INV_X1 g_g8674 (I14816, g8674);
INV_X1 g_I14819 (g8647, I14819);
INV_X1 g_g8675 (I14819, g8675);
INV_X1 g_I14822 (g8649, I14822);
INV_X1 g_g8676 (I14822, g8676);
INV_X1 g_I14825 (g8651, I14825);
INV_X1 g_g8677 (I14825, g8677);
INV_X1 g_I14828 (g8639, I14828);
INV_X1 g_g8678 (I14828, g8678);
INV_X1 g_I14844 (g8641, I14844);
INV_X1 g_g8682 (I14844, g8682);
INV_X1 g_g8683 (g8235, g8683);
INV_X1 g_I14848 (g8625, I14848);
INV_X1 g_g8684 (I14848, g8684);
INV_X1 g_I14851 (g8630, I14851);
INV_X1 g_g8685 (I14851, g8685);
INV_X1 g_I14857 (g8657, I14857);
INV_X1 g_g8689 (I14857, g8689);
INV_X1 g_I14904 (g8629, I14904);
INV_X1 g_g8734 (I14904, g8734);
INV_X1 g_g8743 (g8524, g8743);
INV_X1 g_g8746 (g8524, g8746);
INV_X1 g_g8747 (g8545, g8747);
INV_X1 g_g8750 (g8524, g8750);
INV_X1 g_g8751 (g8545, g8751);
INV_X1 g_g8752 (g8564, g8752);
INV_X1 g_I14925 (g8381, I14925);
INV_X1 g_g8753 (I14925, g8753);
INV_X1 g_g8754 (g8524, g8754);
INV_X1 g_g8755 (g8545, g8755);
INV_X1 g_g8756 (g8564, g8756);
INV_X1 g_g8757 (g8585, g8757);
INV_X1 g_g8759 (g8524, g8759);
INV_X1 g_g8760 (g8545, g8760);
INV_X1 g_g8761 (g8564, g8761);
INV_X1 g_g8762 (g8585, g8762);
INV_X1 g_g8765 (g8524, g8765);
INV_X1 g_g8766 (g8545, g8766);
INV_X1 g_g8767 (g8564, g8767);
INV_X1 g_g8768 (g8585, g8768);
INV_X1 g_g8770 (g8545, g8770);
INV_X1 g_g8771 (g8564, g8771);
INV_X1 g_g8772 (g8585, g8772);
INV_X1 g_I14964 (g8406, I14964);
INV_X1 g_g8774 (I14964, g8774);
INV_X1 g_g8775 (g8564, g8775);
INV_X1 g_g8776 (g8585, g8776);
INV_X1 g_I14974 (g8442, I14974);
INV_X1 g_g8778 (I14974, g8778);
INV_X1 g_g8780 (g8524, g8780);
INV_X1 g_g8781 (g8585, g8781);
INV_X1 g_g8783 (g8524, g8783);
INV_X1 g_g8784 (g8545, g8784);
INV_X1 g_g8786 (g8545, g8786);
INV_X1 g_g8787 (g8564, g8787);
INV_X1 g_g8789 (g8564, g8789);
INV_X1 g_g8790 (g8585, g8790);
INV_X1 g_g8791 (g8585, g8791);
INV_X1 g_I14996 (g8510, I14996);
INV_X1 g_g8792 (I14996, g8792);
INV_X1 g_I15003 (g8633, I15003);
INV_X1 g_g8797 (I15003, g8797);
INV_X1 g_I15007 (g8627, I15007);
INV_X1 g_g8799 (I15007, g8799);
INV_X1 g_I15010 (g8584, I15010);
INV_X1 g_g8800 (I15010, g8800);
INV_X1 g_I15014 (g8607, I15014);
INV_X1 g_g8802 (I15014, g8802);
INV_X1 g_I15062 (g8632, I15062);
INV_X1 g_g8808 (I15062, g8808);
INV_X1 g_I15065 (g8636, I15065);
INV_X1 g_g8809 (I15065, g8809);
INV_X1 g_I15068 (g8638, I15068);
INV_X1 g_g8810 (I15068, g8810);
INV_X1 g_I15160 (g8631, I15160);
INV_X1 g_g8856 (I15160, g8856);
INV_X1 g_I15178 (g8753, I15178);
INV_X1 g_g8864 (I15178, g8864);
INV_X1 g_I15181 (g8734, I15181);
INV_X1 g_g8865 (I15181, g8865);
INV_X1 g_I15184 (g8684, I15184);
INV_X1 g_g8866 (I15184, g8866);
INV_X1 g_I15187 (g8682, I15187);
INV_X1 g_g8867 (I15187, g8867);
INV_X1 g_I15190 (g8685, I15190);
INV_X1 g_g8868 (I15190, g8868);
INV_X1 g_I15193 (g8774, I15193);
INV_X1 g_g8869 (I15193, g8869);
INV_X1 g_I15196 (g8778, I15196);
INV_X1 g_g8870 (I15196, g8870);
INV_X1 g_I15199 (g8792, I15199);
INV_X1 g_g8871 (I15199, g8871);
INV_X1 g_I15202 (g8797, I15202);
INV_X1 g_g8872 (I15202, g8872);
INV_X1 g_I15205 (g8809, I15205);
INV_X1 g_g8873 (I15205, g8873);
INV_X1 g_I15208 (g8810, I15208);
INV_X1 g_g8874 (I15208, g8874);
INV_X1 g_I15211 (g8808, I15211);
INV_X1 g_g8875 (I15211, g8875);
INV_X1 g_I15218 (g8801, I15218);
INV_X1 g_g8880 (I15218, g8880);
INV_X1 g_g8881 (g8683, g8881);
INV_X1 g_I15222 (g8834, I15222);
INV_X1 g_g8882 (I15222, g8882);
INV_X1 g_I15225 (g8689, I15225);
INV_X1 g_g8883 (I15225, g8883);
INV_X1 g_I15308 (g8799, I15308);
INV_X1 g_g8898 (I15308, g8898);
INV_X1 g_I15315 (g8738, I15315);
INV_X1 g_g8903 (I15315, g8903);
INV_X1 g_I15324 (g8779, I15324);
INV_X1 g_g8910 (I15324, g8910);
INV_X1 g_I15329 (g8793, I15329);
INV_X1 g_g8913 (I15329, g8913);
INV_X1 g_I15334 (g8800, I15334);
INV_X1 g_g8916 (I15334, g8916);
INV_X1 g_I15337 (g8802, I15337);
INV_X1 g_g8917 (I15337, g8917);
INV_X1 g_I15340 (g8856, I15340);
INV_X1 g_g8918 (I15340, g8918);
INV_X1 g_I15379 (g8882, I15379);
INV_X1 g_g8955 (I15379, g8955);
INV_X1 g_I15382 (g8883, I15382);
INV_X1 g_g8956 (I15382, g8956);
INV_X1 g_I15385 (g8880, I15385);
INV_X1 g_g8957 (I15385, g8957);
INV_X1 g_I15388 (g8898, I15388);
INV_X1 g_g8958 (I15388, g8958);
INV_X1 g_I15391 (g8917, I15391);
INV_X1 g_g8959 (I15391, g8959);
INV_X1 g_I15394 (g8916, I15394);
INV_X1 g_g8960 (I15394, g8960);
INV_X1 g_I15405 (g8902, I15405);
INV_X1 g_g8967 (I15405, g8967);
INV_X1 g_I15408 (g8896, I15408);
INV_X1 g_g8968 (I15408, g8968);
INV_X1 g_I15411 (g8897, I15411);
INV_X1 g_g8969 (I15411, g8969);
INV_X1 g_I15414 (g8900, I15414);
INV_X1 g_g8970 (I15414, g8970);
INV_X1 g_I15417 (g8893, I15417);
INV_X1 g_g8971 (I15417, g8971);
INV_X1 g_I15420 (g8881, I15420);
INV_X1 g_g8972 (I15420, g8972);
INV_X1 g_I15423 (g8894, I15423);
INV_X1 g_g8973 (I15423, g8973);
INV_X1 g_I15426 (g8895, I15426);
INV_X1 g_g8974 (I15426, g8974);
INV_X1 g_I15429 (g8899, I15429);
INV_X1 g_g8975 (I15429, g8975);
INV_X1 g_I15433 (g8911, I15433);
INV_X1 g_g8977 (I15433, g8977);
INV_X1 g_I15475 (g8901, I15475);
INV_X1 g_g9017 (I15475, g9017);
INV_X1 g_I15478 (g8910, I15478);
INV_X1 g_g9018 (I15478, g9018);
INV_X1 g_I15481 (g8913, I15481);
INV_X1 g_g9019 (I15481, g9019);
INV_X1 g_I15484 (g8918, I15484);
INV_X1 g_g9020 (I15484, g9020);
INV_X1 g_I15492 (g8971, I15492);
INV_X1 g_g9026 (I15492, g9026);
INV_X1 g_I15495 (g8973, I15495);
INV_X1 g_g9027 (I15495, g9027);
INV_X1 g_I15498 (g8974, I15498);
INV_X1 g_g9028 (I15498, g9028);
INV_X1 g_I15501 (g8975, I15501);
INV_X1 g_g9029 (I15501, g9029);
INV_X1 g_I15504 (g8967, I15504);
INV_X1 g_g9030 (I15504, g9030);
INV_X1 g_I15507 (g8968, I15507);
INV_X1 g_g9031 (I15507, g9031);
INV_X1 g_I15510 (g8969, I15510);
INV_X1 g_g9032 (I15510, g9032);
INV_X1 g_I15513 (g8970, I15513);
INV_X1 g_g9033 (I15513, g9033);
INV_X1 g_I15516 (g8977, I15516);
INV_X1 g_g9034 (I15516, g9034);
INV_X1 g_I15519 (g9019, I15519);
INV_X1 g_g9035 (I15519, g9035);
INV_X1 g_I15522 (g9018, I15522);
INV_X1 g_g9036 (I15522, g9036);
INV_X1 g_I15527 (g9020, I15527);
INV_X1 g_g9039 (I15527, g9039);
INV_X1 g_I15530 (g8972, I15530);
INV_X1 g_g9042 (I15530, g9042);
INV_X1 g_I15533 (g9002, I15533);
INV_X1 g_g9043 (I15533, g9043);
INV_X1 g_I15536 (g9004, I15536);
INV_X1 g_g9044 (I15536, g9044);
INV_X1 g_I15539 (g9005, I15539);
INV_X1 g_g9045 (I15539, g9045);
INV_X1 g_I15543 (g9006, I15543);
INV_X1 g_g9047 (I15543, g9047);
INV_X1 g_I15546 (g9007, I15546);
INV_X1 g_g9048 (I15546, g9048);
INV_X1 g_I15550 (g9008, I15550);
INV_X1 g_g9050 (I15550, g9050);
INV_X1 g_I15553 (g9009, I15553);
INV_X1 g_g9051 (I15553, g9051);
INV_X1 g_I15557 (g9010, I15557);
INV_X1 g_g9053 (I15557, g9053);
INV_X1 g_I15562 (g8979, I15562);
INV_X1 g_g9056 (I15562, g9056);
INV_X1 g_I15565 (g8980, I15565);
INV_X1 g_g9057 (I15565, g9057);
INV_X1 g_I15568 (g8981, I15568);
INV_X1 g_g9058 (I15568, g9058);
INV_X1 g_I15571 (g8982, I15571);
INV_X1 g_g9059 (I15571, g9059);
INV_X1 g_I15574 (g8983, I15574);
INV_X1 g_g9060 (I15574, g9060);
INV_X1 g_I15577 (g8984, I15577);
INV_X1 g_g9061 (I15577, g9061);
INV_X1 g_I15580 (g8985, I15580);
INV_X1 g_g9062 (I15580, g9062);
INV_X1 g_I15583 (g8986, I15583);
INV_X1 g_g9063 (I15583, g9063);
INV_X1 g_I15586 (g8987, I15586);
INV_X1 g_g9064 (I15586, g9064);
INV_X1 g_I15589 (g8988, I15589);
INV_X1 g_g9065 (I15589, g9065);
INV_X1 g_I15592 (g8989, I15592);
INV_X1 g_g9066 (I15592, g9066);
INV_X1 g_I15595 (g8990, I15595);
INV_X1 g_g9067 (I15595, g9067);
INV_X1 g_I15598 (g8991, I15598);
INV_X1 g_g9068 (I15598, g9068);
INV_X1 g_I15601 (g8992, I15601);
INV_X1 g_g9069 (I15601, g9069);
INV_X1 g_I15604 (g8993, I15604);
INV_X1 g_g9070 (I15604, g9070);
INV_X1 g_I15607 (g8994, I15607);
INV_X1 g_g9071 (I15607, g9071);
INV_X1 g_I15610 (g8995, I15610);
INV_X1 g_g9072 (I15610, g9072);
INV_X1 g_I15613 (g8996, I15613);
INV_X1 g_g9073 (I15613, g9073);
INV_X1 g_I15616 (g8997, I15616);
INV_X1 g_g9074 (I15616, g9074);
INV_X1 g_I15619 (g8998, I15619);
INV_X1 g_g9075 (I15619, g9075);
INV_X1 g_I15622 (g8999, I15622);
INV_X1 g_g9076 (I15622, g9076);
INV_X1 g_I15625 (g9000, I15625);
INV_X1 g_g9077 (I15625, g9077);
INV_X1 g_I15628 (g9001, I15628);
INV_X1 g_g9078 (I15628, g9078);
INV_X1 g_I15631 (g9003, I15631);
INV_X1 g_g9079 (I15631, g9079);
INV_X1 g_I15635 (g8976, I15635);
INV_X1 g_g9081 (I15635, g9081);
INV_X1 g_I15638 (g8978, I15638);
INV_X1 g_g9082 (I15638, g9082);
INV_X1 g_I15641 (g9017, I15641);
INV_X1 g_g9083 (I15641, g9083);
INV_X1 g_I15645 (g9043, I15645);
INV_X1 g_g9085 (I15645, g9085);
INV_X1 g_I15648 (g9044, I15648);
INV_X1 g_g9086 (I15648, g9086);
INV_X1 g_I15651 (g9056, I15651);
INV_X1 g_g9087 (I15651, g9087);
INV_X1 g_I15654 (g9057, I15654);
INV_X1 g_g9088 (I15654, g9088);
INV_X1 g_I15657 (g9059, I15657);
INV_X1 g_g9089 (I15657, g9089);
INV_X1 g_I15660 (g9062, I15660);
INV_X1 g_g9090 (I15660, g9090);
INV_X1 g_I15663 (g9066, I15663);
INV_X1 g_g9091 (I15663, g9091);
INV_X1 g_I15666 (g9070, I15666);
INV_X1 g_g9092 (I15666, g9092);
INV_X1 g_I15669 (g9045, I15669);
INV_X1 g_g9093 (I15669, g9093);
INV_X1 g_I15672 (g9047, I15672);
INV_X1 g_g9094 (I15672, g9094);
INV_X1 g_I15675 (g9058, I15675);
INV_X1 g_g9095 (I15675, g9095);
INV_X1 g_I15678 (g9060, I15678);
INV_X1 g_g9096 (I15678, g9096);
INV_X1 g_I15681 (g9063, I15681);
INV_X1 g_g9097 (I15681, g9097);
INV_X1 g_I15684 (g9067, I15684);
INV_X1 g_g9098 (I15684, g9098);
INV_X1 g_I15687 (g9071, I15687);
INV_X1 g_g9099 (I15687, g9099);
INV_X1 g_I15690 (g9074, I15690);
INV_X1 g_g9100 (I15690, g9100);
INV_X1 g_I15693 (g9048, I15693);
INV_X1 g_g9101 (I15693, g9101);
INV_X1 g_I15696 (g9050, I15696);
INV_X1 g_g9102 (I15696, g9102);
INV_X1 g_I15699 (g9061, I15699);
INV_X1 g_g9103 (I15699, g9103);
INV_X1 g_I15702 (g9064, I15702);
INV_X1 g_g9104 (I15702, g9104);
INV_X1 g_I15705 (g9068, I15705);
INV_X1 g_g9105 (I15705, g9105);
INV_X1 g_I15708 (g9072, I15708);
INV_X1 g_g9106 (I15708, g9106);
INV_X1 g_I15711 (g9075, I15711);
INV_X1 g_g9107 (I15711, g9107);
INV_X1 g_I15714 (g9077, I15714);
INV_X1 g_g9108 (I15714, g9108);
INV_X1 g_I15717 (g9051, I15717);
INV_X1 g_g9109 (I15717, g9109);
INV_X1 g_I15720 (g9053, I15720);
INV_X1 g_g9110 (I15720, g9110);
INV_X1 g_I15723 (g9065, I15723);
INV_X1 g_g9111 (I15723, g9111);
INV_X1 g_I15726 (g9069, I15726);
INV_X1 g_g9112 (I15726, g9112);
INV_X1 g_I15729 (g9073, I15729);
INV_X1 g_g9113 (I15729, g9113);
INV_X1 g_I15732 (g9076, I15732);
INV_X1 g_g9114 (I15732, g9114);
INV_X1 g_I15735 (g9078, I15735);
INV_X1 g_g9115 (I15735, g9115);
INV_X1 g_I15738 (g9079, I15738);
INV_X1 g_g9116 (I15738, g9116);
INV_X1 g_I15741 (g9083, I15741);
INV_X1 g_g9117 (I15741, g9117);
INV_X1 g_I15747 (g9042, I15747);
INV_X1 g_g9121 (I15747, g9121);
INV_X1 g_I15753 (g9080, I15753);
INV_X1 g_g9125 (I15753, g9125);
INV_X1 g_I15756 (g9081, I15756);
INV_X1 g_g9126 (I15756, g9126);
INV_X1 g_I15759 (g9082, I15759);
INV_X1 g_g9127 (I15759, g9127);
INV_X1 g_I15762 (g9039, I15762);
INV_X1 g_g9128 (I15762, g9128);
INV_X1 g_I15765 (g9039, I15765);
INV_X1 g_g9129 (I15765, g9129);
INV_X1 g_I15770 (g9121, I15770);
INV_X1 g_g9132 (I15770, g9132);
INV_X1 g_I15773 (g9126, I15773);
INV_X1 g_g9133 (I15773, g9133);
INV_X1 g_I15776 (g9127, I15776);
INV_X1 g_g9134 (I15776, g9134);
INV_X1 g_I15784 (g9125, I15784);
INV_X1 g_g9140 (I15784, g9140);
INV_X1 g_g9141 (g9129, g9141);
INV_X1 g_I15791 (g9140, I15791);
INV_X1 g_g9145 (I15791, g9145);
INV_X1 g_g9157 (g9141, g9157);
INV_X1 g_I15803 (g9148, I15803);
INV_X1 g_g9161 (I15803, g9161);
INV_X1 g_I15811 (g9151, I15811);
INV_X1 g_g9177 (I15811, g9177);
INV_X1 g_I15814 (g9154, I15814);
INV_X1 g_g9178 (I15814, g9178);
INV_X1 g_I15824 (g9157, I15824);
INV_X1 g_g9180 (I15824, g9180);
INV_X1 g_g9181 (g9177, g9181);
INV_X1 g_g9182 (g9178, g9182);
INV_X1 g_g9183 (g9161, g9183);
INV_X1 g_I15830 (g9180, I15830);
INV_X1 g_g9184 (I15830, g9184);
INV_X1 g_I15833 (g9162, I15833);
INV_X1 g_g9185 (I15833, g9185);
INV_X1 g_I15836 (g9165, I15836);
INV_X1 g_g9186 (I15836, g9186);
INV_X1 g_I15839 (g9168, I15839);
INV_X1 g_g9187 (I15839, g9187);
INV_X1 g_I15842 (g9171, I15842);
INV_X1 g_g9188 (I15842, g9188);
INV_X1 g_I15845 (g9174, I15845);
INV_X1 g_g9189 (I15845, g9189);
INV_X1 g_g9193 (g9181, g9193);
INV_X1 g_g9194 (g9182, g9194);
INV_X1 g_I15871 (g9184, I15871);
INV_X1 g_g9195 (I15871, g9195);
INV_X1 g_g9196 (g9185, g9196);
INV_X1 g_g9197 (g9186, g9197);
INV_X1 g_g9198 (g9187, g9198);
INV_X1 g_g9199 (g9188, g9199);
INV_X1 g_g9200 (g9189, g9200);
INV_X1 g_g9201 (g9183, g9201);
INV_X1 g_I15894 (g9195, I15894);
INV_X1 g_g9204 (I15894, g9204);
INV_X1 g_g9206 (g9196, g9206);
INV_X1 g_g9207 (g9197, g9207);
INV_X1 g_g9208 (g9198, g9208);
INV_X1 g_g9209 (g9199, g9209);
INV_X1 g_g9210 (g9200, g9210);
INV_X1 g_I15909 (g9201, I15909);
INV_X1 g_g9211 (I15909, g9211);
INV_X1 g_I15912 (g9193, I15912);
INV_X1 g_g9212 (I15912, g9212);
INV_X1 g_I15915 (g9194, I15915);
INV_X1 g_g9213 (I15915, g9213);
INV_X1 g_I15918 (g9211, I15918);
INV_X1 g_g9214 (I15918, g9214);
INV_X1 g_I15921 (g9206, I15921);
INV_X1 g_g9215 (I15921, g9215);
INV_X1 g_I15924 (g9207, I15924);
INV_X1 g_g9216 (I15924, g9216);
INV_X1 g_I15927 (g9208, I15927);
INV_X1 g_g9217 (I15927, g9217);
INV_X1 g_I15930 (g9209, I15930);
INV_X1 g_g9218 (I15930, g9218);
INV_X1 g_I15933 (g9210, I15933);
INV_X1 g_g9219 (I15933, g9219);
INV_X1 g_g9220 (g9205, g9220);
INV_X1 g_I15937 (g9212, I15937);
INV_X1 g_g9221 (I15937, g9221);
INV_X1 g_I15940 (g9213, I15940);
INV_X1 g_g9222 (I15940, g9222);
INV_X1 g_I15943 (g9214, I15943);
INV_X1 g_g9223 (I15943, g9223);
INV_X1 g_I15947 (g9221, I15947);
INV_X1 g_g9227 (I15947, g9227);
INV_X1 g_I15950 (g9222, I15950);
INV_X1 g_g9230 (I15950, g9230);
INV_X1 g_I15953 (g9215, I15953);
INV_X1 g_g9233 (I15953, g9233);
INV_X1 g_I15956 (g9216, I15956);
INV_X1 g_g9234 (I15956, g9234);
INV_X1 g_I15959 (g9217, I15959);
INV_X1 g_g9235 (I15959, g9235);
INV_X1 g_I15962 (g9218, I15962);
INV_X1 g_g9236 (I15962, g9236);
INV_X1 g_I15965 (g9219, I15965);
INV_X1 g_g9237 (I15965, g9237);
INV_X1 g_I15971 (g9233, I15971);
INV_X1 g_g9241 (I15971, g9241);
INV_X1 g_I15974 (g9234, I15974);
INV_X1 g_g9244 (I15974, g9244);
INV_X1 g_I15978 (g9235, I15978);
INV_X1 g_g9248 (I15978, g9248);
INV_X1 g_I15982 (g9236, I15982);
INV_X1 g_g9252 (I15982, g9252);
INV_X1 g_I15985 (g9237, I15985);
INV_X1 g_g9255 (I15985, g9255);
INV_X1 g_I15990 (g9239, I15990);
INV_X1 g_g9260 (I15990, g9260);
INV_X1 g_I16006 (g9261, I16006);
INV_X1 g_g9280 (I16006, g9280);
INV_X1 g_I16009 (g9261, I16009);
INV_X1 g_g9281 (I16009, g9281);
INV_X1 g_I16017 (g9264, I16017);
INV_X1 g_g9297 (I16017, g9297);
INV_X1 g_I16020 (g9264, I16020);
INV_X1 g_g9298 (I16020, g9298);
INV_X1 g_I16023 (g9267, I16023);
INV_X1 g_g9299 (I16023, g9299);
INV_X1 g_I16026 (g9267, I16026);
INV_X1 g_g9300 (I16026, g9300);
INV_X1 g_g9301 (g9260, g9301);
INV_X1 g_g9302 (g9281, g9302);
INV_X1 g_g9303 (g9301, g9303);
INV_X1 g_g9304 (g9298, g9304);
INV_X1 g_I16033 (g9282, I16033);
INV_X1 g_g9305 (I16033, g9305);
INV_X1 g_I16036 (g9282, I16036);
INV_X1 g_g9306 (I16036, g9306);
INV_X1 g_g9307 (g9300, g9307);
INV_X1 g_I16040 (g9285, I16040);
INV_X1 g_g9308 (I16040, g9308);
INV_X1 g_I16043 (g9285, I16043);
INV_X1 g_g9309 (I16043, g9309);
INV_X1 g_I16046 (g9288, I16046);
INV_X1 g_g9310 (I16046, g9310);
INV_X1 g_I16049 (g9288, I16049);
INV_X1 g_g9311 (I16049, g9311);
INV_X1 g_I16052 (g9291, I16052);
INV_X1 g_g9312 (I16052, g9312);
INV_X1 g_I16055 (g9291, I16055);
INV_X1 g_g9313 (I16055, g9313);
INV_X1 g_I16058 (g9294, I16058);
INV_X1 g_g9314 (I16058, g9314);
INV_X1 g_I16061 (g9294, I16061);
INV_X1 g_g9315 (I16061, g9315);
INV_X1 g_g9316 (g9302, g9316);
INV_X1 g_g9317 (g9306, g9317);
INV_X1 g_g9318 (g9304, g9318);
INV_X1 g_g9319 (g9309, g9319);
INV_X1 g_g9320 (g9307, g9320);
INV_X1 g_g9321 (g9311, g9321);
INV_X1 g_g9322 (g9313, g9322);
INV_X1 g_g9323 (g9315, g9323);
INV_X1 g_I16072 (g9303, I16072);
INV_X1 g_g9324 (I16072, g9324);
INV_X1 g_g9329 (g9317, g9329);
INV_X1 g_g9330 (g9319, g9330);
INV_X1 g_g9331 (g9321, g9331);
INV_X1 g_g9332 (g9322, g9332);
INV_X1 g_g9333 (g9323, g9333);
INV_X1 g_I16084 (g9324, I16084);
INV_X1 g_g9336 (I16084, g9336);
INV_X1 g_I16090 (g9336, I16090);
INV_X1 g_g9340 (I16090, g9340);
INV_X1 g_I16100 (g9338, I16100);
INV_X1 g_g9350 (I16100, g9350);
INV_X1 g_I16103 (g9339, I16103);
INV_X1 g_g9351 (I16103, g9351);
INV_X1 g_I16107 (g9337, I16107);
INV_X1 g_g9353 (I16107, g9353);
INV_X1 g_I16116 (g9350, I16116);
INV_X1 g_g9360 (I16116, g9360);
INV_X1 g_I16119 (g9351, I16119);
INV_X1 g_g9361 (I16119, g9361);
INV_X1 g_I16122 (g9353, I16122);
INV_X1 g_g9362 (I16122, g9362);
INV_X1 g_I16126 (g9354, I16126);
INV_X1 g_g9366 (I16126, g9366);
INV_X1 g_I16129 (g9355, I16129);
INV_X1 g_g9367 (I16129, g9367);
INV_X1 g_I16132 (g9356, I16132);
INV_X1 g_g9368 (I16132, g9368);
INV_X1 g_I16135 (g9357, I16135);
INV_X1 g_g9369 (I16135, g9369);
INV_X1 g_I16138 (g9358, I16138);
INV_X1 g_g9370 (I16138, g9370);
INV_X1 g_I16142 (g9366, I16142);
INV_X1 g_g9372 (I16142, g9372);
INV_X1 g_I16145 (g9367, I16145);
INV_X1 g_g9373 (I16145, g9373);
INV_X1 g_I16148 (g9368, I16148);
INV_X1 g_g9374 (I16148, g9374);
INV_X1 g_I16151 (g9369, I16151);
INV_X1 g_g9375 (I16151, g9375);
INV_X1 g_I16154 (g9370, I16154);
INV_X1 g_g9376 (I16154, g9376);
INV_X1 g_I16158 (g9363, I16158);
INV_X1 g_g9378 (I16158, g9378);
INV_X1 g_I16161 (g9363, I16161);
INV_X1 g_g9379 (I16161, g9379);
INV_X1 g_g9380 (g9379, g9380);
INV_X1 g_I16165 (g9377, I16165);
INV_X1 g_g9381 (I16165, g9381);
INV_X1 g_I16168 (g9381, I16168);
INV_X1 g_g9382 (I16168, g9382);
INV_X1 g_g9383 (g9380, g9383);
INV_X1 g_I16173 (g9382, I16173);
INV_X1 g_g9385 (I16173, g9385);
INV_X1 g_I16176 (g9385, I16176);
INV_X1 g_g9386 (I16176, g9386);
INV_X1 g_I16180 (g9387, I16180);
INV_X1 g_g9388 (I16180, g9388);
INV_X1 g_I16183 (g9388, I16183);
INV_X1 g_g9389 (I16183, g9389);
AND2_X1 g_g1714 (g1454, g1450, g1714);
AND2_X1 g_g1725 (g1409, g1416, g1725);
AND2_X1 g_g1728 (g1432, g1439, g1728);
AND2_X1 g_g1733 (g1489, g1481, g1733);
AND2_X1 g_g1739 (g803, g799, g1739);
AND2_X1 g_g1753 (g819, g815, g1753);
AND2_X1 g_g1834 (g933, g929, g1834);
AND2_X1 g_g1844 (g792, g795, g1844);
AND2_X1 g_g1898 (g959, g955, g1898);
AND2_X1 g_g1913 (g1528, g1532, g1913);
AND2_X1 g_g1919 (g1098, g1087, g1919);
AND2_X1 g_g2386 (g1130, g1092, g2386);
AND2_X1 g_g2768 (g1597, g973, g2768);
AND2_X1 g_g2781 (g1600, g976, g2781);
AND2_X1 g_g2827 (g1889, g1690, g2827);
AND2_X1 g_g2889 (g1612, g1077, g2889);
AND2_X1 g_g2912 (g1080, g1945, g2912);
AND2_X1 g_g2935 (g1612, g1077, g2935);
AND2_X1 g_g2949 (g822, g1753, g2949);
AND2_X1 g_g2952 (g2474, g2215, g2952);
AND2_X1 g_g2972 (g2397, g2407, g2972);
AND2_X1 g_g2979 (g1494, g1733, g2979);
AND2_X1 g_g2986 (g806, g1739, g2986);
AND2_X1 g_g3002 (g871, g1834, g3002);
AND2_X1 g_g3049 (g2274, g1844, g3049);
AND2_X1 g_g3081 (g1682, g1616, g3081);
AND2_X1 g_g3094 (g945, g1898, g3094);
AND2_X1 g_g3188 (g2298, g2316, g3188);
AND2_X1 g_g3190 (g1658, g2424, g3190);
AND2_X1 g_g3222 (g1537, g1913, g3222);
AND2_X1 g_g3226 (g1102, g1919, g3226);
AND2_X1 g_g3229 (g1728, g2015, g3229);
AND4_X1 g_g3258 (g2298, g2316, g2334, g2354, g3258);
AND2_X1 g_g3259 (g1976, g1960, g3259);
AND3_X1 g_g3313 (g2334, g2316, g2298, g3313);
AND3_X1 g_g3429 (g1454, g1838, g1444, g3429);
AND2_X1 g_g3466 (g936, g2557, g3466);
AND2_X1 g_g3509 (g1637, g1616, g3509);
AND2_X1 g_g3614 (g1134, g2386, g3614);
AND2_X1 g_g3984 (g2403, g3085, g3984);
AND2_X1 g_g4038 (g825, g2949, g4038);
AND2_X1 g_g4047 (g1272, g3503, g4047);
AND2_X1 g_g4048 (g1288, g3513, g4048);
AND2_X1 g_g4049 (g141, g3514, g4049);
AND2_X1 g_g4052 (g1276, g3522, g4052);
AND2_X1 g_g4053 (g1292, g3523, g4053);
AND2_X1 g_g4054 (g3767, g2424, g4054);
AND2_X1 g_g4058 (g3656, g2407, g4058);
AND2_X1 g_g4059 (g1499, g2979, g4059);
AND2_X1 g_g4062 (g809, g2986, g4062);
AND2_X1 g_g4066 (g1280, g3532, g4066);
AND2_X1 g_g4067 (g133, g3539, g4067);
AND2_X1 g_g4068 (g121, g3540, g4068);
AND2_X1 g_g4073 (g1300, g3567, g4073);
AND2_X1 g_g4074 (g137, g3573, g4074);
AND2_X1 g_g4077 (g1284, g3582, g4077);
AND4_X1 g_g4078 (g3753, g3732, g3712, g3700, g4078);
AND2_X1 g_g4082 (g1296, g3604, g4082);
AND2_X1 g_g4083 (g125, g3610, g4083);
AND2_X1 g_g4086 (g103, g3629, g4086);
AND2_X1 g_g4091 (g129, g3639, g4091);
AND2_X1 g_g4097 (g2624, g2614, g4097);
AND2_X1 g_g4098 (g985, g3790, g4098);
AND2_X1 g_g4099 (g117, g3647, g4099);
AND2_X1 g_g4100 (g113, g3648, g4100);
AND2_X1 g_g4101 (g108, g3649, g4101);
AND2_X1 g_g4107 (g2625, g2615, g4107);
AND2_X1 g_g4108 (g782, g3655, g4108);
AND2_X1 g_g4109 (g990, g3790, g4109);
AND2_X1 g_g4117 (g2626, g2616, g4117);
AND2_X1 g_g4118 (g995, g3790, g4118);
AND2_X1 g_g4123 (g2627, g2617, g4123);
AND2_X1 g_g4124 (g2641, g2640, g4124);
AND2_X1 g_g4127 (g2628, g2618, g4127);
AND2_X1 g_g4128 (g98, g3693, g4128);
AND2_X1 g_g4129 (g2629, g2621, g4129);
AND2_X1 g_g4131 (g2630, g2622, g4131);
AND2_X1 g_g4132 (g2637, g2633, g4132);
AND2_X1 g_g4133 (g2631, g2623, g4133);
AND4_X1 g_I7994 (g3430, g3398, g3359, g3341, I7994);
AND4_X1 g_I7995 (g2074, g3287, g2020, g3238, I7995);
AND2_X1 g_g4135 (I7994, I7995, g4135);
AND2_X1 g_g4138 (g2638, g2634, g4138);
AND4_X1 g_I8000 (g3430, g3398, g3359, g3341, I8000);
AND4_X1 g_I8001 (g2074, g3287, g2020, g1987, I8001);
AND2_X1 g_g4139 (I8000, I8001, g4139);
AND4_X1 g_I8005 (g3430, g3398, g3359, g2106, I8005);
AND4_X1 g_I8006 (g2074, g3287, g2020, g3238, I8006);
AND2_X1 g_g4142 (I8005, I8006, g4142);
AND2_X1 g_g4145 (g2639, g2635, g4145);
AND4_X1 g_I8014 (g3430, g3398, g3359, g3341, I8014);
AND4_X1 g_I8015 (g2074, g2057, g3264, g3238, I8015);
AND2_X1 g_g4147 (I8014, I8015, g4147);
AND4_X1 g_I8019 (g3430, g3398, g3359, g2106, I8019);
AND4_X1 g_I8020 (g2074, g3287, g2020, g1987, I8020);
AND2_X1 g_g4150 (I8019, I8020, g4150);
AND2_X1 g_g4154 (g1098, g3495, g4154);
AND4_X1 g_I8028 (g3430, g3398, g3359, g3341, I8028);
AND4_X1 g_I8029 (g2074, g2057, g3264, g1987, I8029);
AND2_X1 g_g4155 (I8028, I8029, g4155);
AND4_X1 g_I8033 (g3430, g3398, g3359, g2106, I8033);
AND4_X1 g_I8034 (g2074, g2057, g3264, g3238, I8034);
AND2_X1 g_g4158 (I8033, I8034, g4158);
AND2_X1 g_g4159 (g1102, g3498, g4159);
AND4_X1 g_I8040 (g3430, g3398, g3359, g3341, I8040);
AND4_X1 g_I8041 (g2074, g2057, g2020, g3238, I8041);
AND2_X1 g_g4163 (I8040, I8041, g4163);
AND4_X1 g_I8045 (g3430, g3398, g3359, g2106, I8045);
AND4_X1 g_I8046 (g2074, g2057, g3264, g1987, I8046);
AND2_X1 g_g4166 (I8045, I8046, g4166);
AND2_X1 g_g4167 (g2783, g1616, g4167);
AND2_X1 g_g4168 (g1106, g3500, g4168);
AND4_X1 g_I8052 (g2162, g2149, g2137, g2106, I8052);
AND4_X1 g_I8053 (g3316, g3287, g3264, g3238, I8053);
AND2_X1 g_g4169 (I8052, I8053, g4169);
AND4_X1 g_I8057 (g3430, g3398, g3359, g3341, I8057);
AND4_X1 g_I8058 (g2074, g2057, g2020, g1987, I8058);
AND2_X1 g_g4172 (I8057, I8058, g4172);
AND2_X1 g_g4175 (g1110, g3502, g4175);
AND4_X1 g_I8063 (g2162, g2149, g2137, g2106, I8063);
AND4_X1 g_I8064 (g3316, g3287, g3264, g1987, I8064);
AND2_X1 g_g4176 (I8063, I8064, g4176);
AND2_X1 g_g4180 (g1114, g3511, g4180);
AND2_X1 g_g4181 (g1142, g3512, g4181);
AND4_X1 g_I8071 (g2162, g2149, g2137, g2106, I8071);
AND4_X1 g_I8072 (g3316, g3287, g2020, g3238, I8072);
AND2_X1 g_g4182 (I8071, I8072, g4182);
AND2_X1 g_g4185 (g2636, g2632, g4185);
AND2_X1 g_g4186 (g1118, g3520, g4186);
AND4_X1 g_I8078 (g2162, g2149, g2137, g2106, I8078);
AND4_X1 g_I8079 (g3316, g3287, g2020, g1987, I8079);
AND2_X1 g_g4187 (I8078, I8079, g4187);
AND2_X1 g_g4190 (g1122, g3527, g4190);
AND2_X1 g_g4192 (g1126, g3531, g4192);
AND2_X1 g_g4193 (g145, g2727, g4193);
AND4_X1 g_I8089 (g2162, g2149, g2137, g2106, I8089);
AND4_X1 g_I8090 (g3316, g2057, g2020, g3238, I8090);
AND2_X1 g_g4194 (I8089, I8090, g4194);
AND2_X1 g_g4199 (g93, g2769, g4199);
AND4_X1 g_I8108 (g2162, g2149, g2137, g2106, I8108);
AND4_X1 g_I8109 (g2074, g3287, g3264, g3238, I8109);
AND2_X1 g_g4201 (I8108, I8109, g4201);
AND4_X1 g_I8114 (g2162, g2149, g2137, g2106, I8114);
AND4_X1 g_I8115 (g2074, g3287, g3264, g1987, I8115);
AND2_X1 g_g4216 (I8114, I8115, g4216);
AND4_X1 g_g4220 (g3533, g3549, g3568, g3583, g4220);
AND3_X1 g_I8127 (g2699, g2674, g2677, I8127);
AND3_X1 g_g4224 (g2680, g2683, I8127, g4224);
AND4_X1 g_g4225 (g2686, g2689, g2692, g2695, g4225);
AND3_X1 g_I8143 (g2674, g2677, g2680, I8143);
AND3_X1 g_g4230 (g2683, g3491, I8143, g4230);
AND2_X1 g_g4236 (g3260, g3221, g4236);
AND3_X1 g_I8157 (g2686, g2689, g2692, I8157);
AND3_X1 g_g4238 (g2695, g2698, I8157, g4238);
AND2_X1 g_g4239 (g1541, g3222, g4239);
AND2_X1 g_g4246 (g1106, g3226, g4246);
AND3_X1 g_g4254 (g3583, g3568, g3549, g4254);
AND4_X1 g_I8186 (g3778, g3549, g3568, g3583, I8186);
AND4_X1 g_g4255 (g3605, g3644, g3635, I8186, g4255);
AND2_X1 g_g4268 (g2216, g2655, g4268);
AND3_X1 g_I8209 (g2298, g2316, g2334, I8209);
AND3_X1 g_g4269 (g2354, g3563, I8209, g4269);
AND2_X1 g_g4271 (g3666, g3684, g4271);
AND2_X1 g_g4272 (g3233, g3286, g4272);
AND2_X1 g_g4276 (g2216, g2618, g4276);
AND2_X1 g_g4282 (g3549, g3568, g4282);
AND2_X1 g_g4284 (g3260, g3314, g4284);
AND3_X1 g_I8237 (g2298, g2316, g2354, I8237);
AND4_X1 g_g4287 (g3563, g2334, g3579, I8237, g4287);
AND4_X1 g_I8240 (g2298, g2316, g2334, g2354, I8240);
AND4_X1 g_g4288 (g3563, g3579, g3603, I8240, g4288);
AND2_X1 g_g4299 (g3233, g3358, g4299);
AND3_X1 g_g4302 (g3086, g3659, g3124, g4302);
AND2_X1 g_g4304 (g2784, g3779, g4304);
AND4_X1 g_g4312 (g3666, g3684, g3694, g3707, g4312);
AND3_X1 g_g4314 (g3694, g3684, g3666, g4314);
AND3_X1 g_I8288 (g3666, g3684, g3694, I8288);
AND3_X1 g_g4315 (g3707, g3728, I8288, g4315);
AND4_X1 g_g4317 (g878, g3086, g1857, g3659, g4317);
AND3_X1 g_I8296 (g3666, g3684, g3707, I8296);
AND4_X1 g_g4319 (g3728, g3694, g3750, I8296, g4319);
AND4_X1 g_I8299 (g3666, g3684, g3694, g3707, I8299);
AND4_X1 g_g4320 (g3728, g3750, g3768, I8299, g4320);
AND2_X1 g_g4327 (g2959, g1867, g4327);
AND2_X1 g_g4333 (g1087, g2782, g4333);
AND2_X1 g_g4334 (g225, g3097, g4334);
AND2_X1 g_g4342 (g228, g3097, g4342);
AND2_X1 g_g4343 (g306, g3131, g4343);
AND2_X1 g_g4351 (g309, g3131, g4351);
AND2_X1 g_g4352 (g387, g3160, g4352);
AND2_X1 g_g4355 (g390, g3160, g4355);
AND2_X1 g_g4356 (g468, g3192, g4356);
AND2_X1 g_g4361 (g471, g3192, g4361);
AND2_X1 g_g4365 (g237, g3097, g4365);
AND2_X1 g_g4366 (g216, g3097, g4366);
AND2_X1 g_g4367 (g240, g3097, g4367);
AND2_X1 g_g4368 (g318, g3131, g4368);
AND2_X1 g_g4369 (g580, g2845, g4369);
AND2_X1 g_g4375 (g219, g3097, g4375);
AND2_X1 g_g4376 (g243, g3097, g4376);
AND2_X1 g_g4377 (g297, g3131, g4377);
AND2_X1 g_g4378 (g321, g3131, g4378);
AND2_X1 g_g4379 (g399, g3160, g4379);
AND2_X1 g_g4380 (g584, g2845, g4380);
AND2_X1 g_g4383 (g222, g3097, g4383);
AND2_X1 g_g4384 (g246, g3097, g4384);
AND2_X1 g_g4385 (g300, g3131, g4385);
AND2_X1 g_g4386 (g324, g3131, g4386);
AND2_X1 g_g4387 (g378, g3160, g4387);
AND2_X1 g_g4388 (g402, g3160, g4388);
AND2_X1 g_g4389 (g480, g3192, g4389);
AND2_X1 g_g4390 (g560, g2845, g4390);
AND2_X1 g_g4391 (g249, g3097, g4391);
AND2_X1 g_g4392 (g303, g3131, g4392);
AND2_X1 g_g4393 (g327, g3131, g4393);
AND2_X1 g_g4394 (g381, g3160, g4394);
AND2_X1 g_g4395 (g405, g3160, g4395);
AND2_X1 g_g4396 (g459, g3192, g4396);
AND2_X1 g_g4397 (g483, g3192, g4397);
AND2_X1 g_g4398 (g567, g2845, g4398);
AND2_X1 g_g4400 (g1138, g3614, g4400);
AND4_X1 g_I8400 (g3430, g3398, g3359, g3341, I8400);
AND4_X1 g_I8401 (g3316, g3287, g3264, g3238, I8401);
AND2_X1 g_g4403 (I8400, I8401, g4403);
AND2_X1 g_g4407 (g252, g3097, g4407);
AND2_X1 g_g4408 (g330, g3131, g4408);
AND2_X1 g_g4409 (g384, g3160, g4409);
AND2_X1 g_g4410 (g408, g3160, g4410);
AND2_X1 g_g4411 (g462, g3192, g4411);
AND2_X1 g_g4412 (g486, g3192, g4412);
AND4_X1 g_I8412 (g3430, g3398, g3359, g3341, I8412);
AND4_X1 g_I8413 (g3316, g3287, g3264, g1987, I8413);
AND2_X1 g_g4414 (I8412, I8413, g4414);
AND4_X1 g_I8417 (g3430, g3398, g3359, g2106, I8417);
AND4_X1 g_I8418 (g3316, g3287, g3264, g3238, I8418);
AND2_X1 g_g4417 (I8417, I8418, g4417);
AND2_X1 g_g4420 (g275, g3097, g4420);
AND2_X1 g_g4421 (g333, g3131, g4421);
AND2_X1 g_g4422 (g411, g3160, g4422);
AND2_X1 g_g4423 (g465, g3192, g4423);
AND2_X1 g_g4424 (g489, g3192, g4424);
AND2_X1 g_g4425 (g536, g2845, g4425);
AND4_X1 g_I8431 (g3430, g3398, g3359, g3341, I8431);
AND4_X1 g_I8432 (g3316, g3287, g2020, g3238, I8432);
AND2_X1 g_g4427 (I8431, I8432, g4427);
AND4_X1 g_I8436 (g3430, g3398, g3359, g2106, I8436);
AND4_X1 g_I8437 (g3316, g3287, g3264, g1987, I8437);
AND2_X1 g_g4430 (I8436, I8437, g4430);
AND2_X1 g_g4433 (g278, g3097, g4433);
AND2_X1 g_g4434 (g356, g3131, g4434);
AND2_X1 g_g4435 (g414, g3160, g4435);
AND2_X1 g_g4436 (g492, g3192, g4436);
AND2_X1 g_g4437 (g540, g2845, g4437);
AND4_X1 g_I8455 (g3430, g3398, g3359, g3341, I8455);
AND4_X1 g_I8456 (g3316, g3287, g2020, g1987, I8456);
AND2_X1 g_g4445 (I8455, I8456, g4445);
AND4_X1 g_I8460 (g3430, g3398, g3359, g2106, I8460);
AND4_X1 g_I8461 (g3316, g3287, g2020, g3238, I8461);
AND2_X1 g_g4448 (I8460, I8461, g4448);
AND2_X1 g_g4451 (g359, g3131, g4451);
AND2_X1 g_g4452 (g437, g3160, g4452);
AND2_X1 g_g4453 (g495, g3192, g4453);
AND2_X1 g_g4454 (g544, g2845, g4454);
AND4_X1 g_I8490 (g3430, g3398, g3359, g3341, I8490);
AND4_X1 g_I8491 (g3316, g2057, g3264, g3238, I8491);
AND2_X1 g_g4466 (I8490, I8491, g4466);
AND4_X1 g_I8495 (g3430, g3398, g3359, g2106, I8495);
AND4_X1 g_I8496 (g3316, g3287, g2020, g1987, I8496);
AND2_X1 g_g4469 (I8495, I8496, g4469);
AND2_X1 g_g4472 (g440, g3160, g4472);
AND2_X1 g_g4473 (g518, g3192, g4473);
AND4_X1 g_I8523 (g3430, g3398, g3359, g3341, I8523);
AND4_X1 g_I8524 (g3316, g2057, g3264, g1987, I8524);
AND2_X1 g_g4483 (I8523, I8524, g4483);
AND4_X1 g_I8528 (g3430, g3398, g3359, g2106, I8528);
AND4_X1 g_I8529 (g3316, g2057, g3264, g3238, I8529);
AND2_X1 g_g4486 (I8528, I8529, g4486);
AND2_X1 g_g4490 (g521, g3192, g4490);
AND2_X1 g_g4491 (g557, g2845, g4491);
AND4_X1 g_I8546 (g3430, g3398, g3359, g3341, I8546);
AND4_X1 g_I8547 (g3316, g2057, g2020, g3238, I8547);
AND2_X1 g_g4494 (I8546, I8547, g4494);
AND4_X1 g_I8551 (g3430, g3398, g3359, g2106, I8551);
AND4_X1 g_I8552 (g3316, g2057, g3264, g1987, I8552);
AND2_X1 g_g4497 (I8551, I8552, g4497);
AND4_X1 g_I8568 (g3430, g3398, g3359, g3341, I8568);
AND4_X1 g_I8569 (g3316, g2057, g2020, g1987, I8569);
AND2_X1 g_g4504 (I8568, I8569, g4504);
AND4_X1 g_I8573 (g3430, g3398, g3359, g2106, I8573);
AND4_X1 g_I8574 (g3316, g2057, g2020, g3238, I8574);
AND2_X1 g_g4507 (I8573, I8574, g4507);
AND4_X1 g_I8588 (g3430, g3398, g3359, g3341, I8588);
AND4_X1 g_I8589 (g2074, g3287, g3264, g3238, I8589);
AND2_X1 g_g4514 (I8588, I8589, g4514);
AND4_X1 g_I8593 (g3430, g3398, g3359, g2106, I8593);
AND4_X1 g_I8594 (g3316, g2057, g2020, g1987, I8594);
AND2_X1 g_g4517 (I8593, I8594, g4517);
AND2_X1 g_g4526 (g2642, g741, g4526);
AND4_X1 g_I8612 (g3430, g3398, g3359, g3341, I8612);
AND4_X1 g_I8613 (g2074, g3287, g3264, g1987, I8613);
AND2_X1 g_g4529 (I8612, I8613, g4529);
AND4_X1 g_I8617 (g3430, g3398, g3359, g2106, I8617);
AND4_X1 g_I8618 (g2074, g3287, g3264, g3238, I8618);
AND2_X1 g_g4532 (I8617, I8618, g4532);
AND2_X1 g_g4546 (g2643, g746, g4546);
AND4_X1 g_I8642 (g3430, g3398, g3359, g2106, I8642);
AND4_X1 g_I8643 (g2074, g3287, g3264, g1987, I8643);
AND2_X1 g_g4549 (I8642, I8643, g4549);
AND2_X1 g_g4681 (g4255, g3533, g4681);
AND2_X1 g_g4690 (g4081, g3078, g4690);
AND2_X1 g_g4691 (g4219, g1690, g4691);
AND2_X1 g_g4699 (g1557, g4276, g4699);
AND2_X1 g_g4702 (g4243, g1690, g4702);
AND2_X1 g_g4705 (g190, g3986, g4705);
AND2_X1 g_g4707 (g812, g4062, g4707);
AND2_X1 g_g4711 (g190, g4072, g4711);
AND2_X1 g_g4712 (g1179, g4276, g4712);
AND2_X1 g_g4720 (g190, g4055, g4720);
AND2_X1 g_g4724 (g828, g4038, g4724);
AND2_X1 g_g4728 (g190, g4179, g4728);
AND2_X1 g_g4729 (g1504, g4059, g4729);
AND2_X1 g_g4740 (g2242, g4275, g4740);
AND2_X1 g_g4743 (g3518, g4286, g4743);
AND2_X1 g_g4744 (g3525, g4296, g4744);
AND2_X1 g_g4778 (g4169, g1760, g4778);
AND2_X1 g_g4779 (g4176, g1760, g4779);
AND2_X1 g_g4781 (g4182, g1760, g4781);
AND2_X1 g_g4782 (g4187, g1760, g4782);
AND2_X1 g_g4783 (g948, g4527, g4783);
AND2_X1 g_g4785 (g1678, g4202, g4785);
AND2_X1 g_g4787 (g953, g4547, g4787);
AND2_X1 g_g4789 (g2751, g4202, g4789);
AND2_X1 g_g4791 (g949, g4562, g4791);
AND2_X1 g_g4793 (g3887, g4202, g4793);
AND2_X1 g_g4794 (g954, g4574, g4794);
AND2_X1 g_g4796 (g950, g4584, g4796);
AND2_X1 g_g4797 (g3893, g1616, g4797);
AND2_X1 g_g4798 (g4216, g1760, g4798);
AND2_X1 g_g4799 (g951, g4596, g4799);
AND2_X1 g_g4804 (g952, g3876, g4804);
AND2_X1 g_g4814 (g150, g4265, g4814);
AND3_X1 g_I9166 (g4041, g2595, g2584, I9166);
AND3_X1 g_g4819 (g2573, g2562, I9166, g4819);
AND3_X1 g_g4823 (g4238, g4230, g174, g4823);
AND2_X1 g_g4825 (g4228, g1964, g4825);
AND2_X1 g_g4826 (g1545, g4239, g4826);
AND2_X1 g_g4830 (g4288, g3723, g4830);
AND2_X1 g_g4832 (g1110, g4246, g4832);
AND3_X1 g_I9202 (g2605, g4044, g2584, I9202);
AND3_X1 g_g4837 (g2573, g2562, I9202, g4837);
AND2_X1 g_g4838 (g4517, g1760, g4838);
AND2_X1 g_g4840 (g4235, g1980, g4840);
AND2_X1 g_g4868 (g4227, g4160, g4868);
AND3_X1 g_g4872 (g1924, g4225, g4224, g4872);
AND4_X1 g_g4877 (g3746, g3723, g4288, g3764, g4877);
AND3_X1 g_I9222 (g4041, g4044, g2584, I9222);
AND3_X1 g_g4878 (g2573, g2562, I9222, g4878);
AND3_X1 g_g4883 (g3746, g3723, g4288, g4883);
AND3_X1 g_I9261 (g3777, g3764, g3746, I9261);
AND3_X1 g_g4901 (g3723, g4288, I9261, g4901);
AND4_X1 g_g4902 (g4304, g2770, g2746, g2728, g4902);
AND2_X1 g_g4906 (g4320, g2728, g4906);
AND4_X1 g_g4933 (g2746, g2728, g4320, g2770, g4933);
AND2_X1 g_g4936 (g214, g3888, g4936);
AND2_X1 g_g4937 (g3086, g4309, g4937);
AND2_X1 g_g4955 (g215, g3891, g4955);
AND2_X1 g_g4956 (g295, g3892, g4956);
AND3_X1 g_g4957 (g2746, g2728, g4320, g4957);
AND2_X1 g_g4958 (g296, g3897, g4958);
AND2_X1 g_g4959 (g376, g3898, g4959);
AND2_X1 g_g4961 (g377, g3904, g4961);
AND2_X1 g_g4962 (g457, g3905, g4962);
AND2_X1 g_g4968 (g4403, g1760, g4968);
AND2_X1 g_g4969 (g4362, g2216, g4969);
AND2_X1 g_g5001 (g458, g3912, g5001);
AND3_X1 g_I9330 (g2784, g2770, g2746, I9330);
AND3_X1 g_g5005 (g2728, g4320, I9330, g5005);
AND2_X1 g_g5008 (g231, g3920, g5008);
AND2_X1 g_g5017 (g211, g3928, g5017);
AND2_X1 g_g5018 (g232, g3930, g5018);
AND2_X1 g_g5019 (g312, g3933, g5019);
AND2_X1 g_g5020 (g579, g3937, g5020);
AND2_X1 g_g5029 (g212, g3945, g5029);
AND2_X1 g_g5030 (g233, g3946, g5030);
AND2_X1 g_g5031 (g292, g3948, g5031);
AND2_X1 g_g5032 (g313, g3950, g5032);
AND2_X1 g_g5033 (g393, g3953, g5033);
AND2_X1 g_g5034 (g583, g3956, g5034);
AND2_X1 g_g5043 (g213, g3958, g5043);
AND2_X1 g_g5044 (g234, g3959, g5044);
AND2_X1 g_g5045 (g293, g3961, g5045);
AND2_X1 g_g5046 (g314, g3962, g5046);
AND2_X1 g_g5047 (g373, g3964, g5047);
AND2_X1 g_g5048 (g394, g3966, g5048);
AND2_X1 g_g5049 (g474, g3969, g5049);
AND2_X1 g_g5050 (g587, g3970, g5050);
AND2_X1 g_g5062 (g235, g3973, g5062);
AND2_X1 g_g5063 (g294, g3974, g5063);
AND2_X1 g_g5064 (g315, g3975, g5064);
AND2_X1 g_g5065 (g374, g3977, g5065);
AND2_X1 g_g5066 (g395, g3978, g5066);
AND2_X1 g_g5067 (g454, g3980, g5067);
AND2_X1 g_g5068 (g475, g3982, g5068);
AND2_X1 g_g5069 (g566, g3983, g5069);
AND2_X1 g_g5077 (g236, g3988, g5077);
AND2_X1 g_g5078 (g316, g3989, g5078);
AND2_X1 g_g5079 (g375, g3990, g5079);
AND2_X1 g_g5080 (g396, g3991, g5080);
AND2_X1 g_g5081 (g455, g3993, g5081);
AND2_X1 g_g5082 (g476, g3994, g5082);
AND2_X1 g_g5089 (g273, g3998, g5089);
AND2_X1 g_g5090 (g317, g4000, g5090);
AND2_X1 g_g5091 (g397, g4001, g5091);
AND2_X1 g_g5092 (g456, g4002, g5092);
AND2_X1 g_g5093 (g477, g4003, g5093);
AND2_X1 g_g5094 (g535, g4004, g5094);
AND2_X1 g_g5096 (g1149, g4400, g5096);
AND2_X1 g_g5104 (g274, g4010, g5104);
AND2_X1 g_g5105 (g354, g4013, g5105);
AND2_X1 g_g5106 (g398, g4015, g5106);
AND2_X1 g_g5107 (g478, g4016, g5107);
AND2_X1 g_g5108 (g539, g4017, g5108);
AND2_X1 g_g5116 (g355, g4021, g5116);
AND2_X1 g_g5117 (g435, g4024, g5117);
AND2_X1 g_g5118 (g479, g4026, g5118);
AND2_X1 g_g5119 (g543, g4027, g5119);
AND2_X1 g_g5122 (g436, g4030, g5122);
AND2_X1 g_g5123 (g516, g4033, g5123);
AND2_X1 g_g5125 (g517, g4036, g5125);
AND2_X1 g_g5126 (g556, g4037, g5126);
AND4_X1 g_I9534 (g3019, g3029, g3038, g3052, I9534);
AND4_X1 g_I9535 (g3062, g2712, g4253, g2752, I9535);
AND2_X1 g_g5132 (I9534, I9535, g5132);
AND2_X1 g_g5142 (g1677, g4202, g5142);
AND2_X1 g_g5287 (g786, g4724, g5287);
AND2_X1 g_g5298 (g1912, g4814, g5298);
AND2_X1 g_g5313 (g4820, g2407, g5313);
AND2_X1 g_g5314 (g1509, g4729, g5314);
AND2_X1 g_g5334 (g4887, g2424, g5334);
AND2_X1 g_g5425 (g1528, g4916, g5425);
AND2_X1 g_g5428 (g775, g4707, g5428);
AND2_X1 g_g5432 (g1537, g4921, g5432);
AND2_X1 g_g5436 (g1541, g4926, g5436);
AND2_X1 g_g5438 (g1545, g4932, g5438);
AND2_X1 g_g5441 (g4870, g3497, g5441);
AND2_X1 g_g5442 (g4679, g4202, g5442);
AND2_X1 g_g5443 (g1549, g4935, g5443);
AND2_X1 g_g5452 (g4876, g3499, g5452);
AND2_X1 g_g5458 (g4686, g1616, g5458);
AND2_X1 g_g5475 (g3801, g5022, g5475);
AND2_X1 g_g5479 (g5141, g5037, g5479);
AND2_X1 g_g5484 (g1037, g5096, g5484);
AND2_X1 g_g5489 (g4912, g5053, g5489);
AND2_X1 g_g5513 (g4889, g5071, g5513);
AND2_X1 g_g5547 (g4814, g1819, g5547);
AND2_X1 g_g5548 (g1549, g4826, g5548);
AND2_X1 g_g5552 (g1114, g4832, g5552);
AND2_X1 g_g5560 (g3390, g5036, g5560);
AND2_X1 g_g5563 (g3390, g5070, g5563);
AND2_X1 g_g5570 (g1759, g4841, g5570);
AND2_X1 g_g5573 (g3011, g4841, g5573);
AND2_X1 g_g5579 (g4090, g4841, g5579);
AND2_X1 g_g5583 (g1775, g4969, g5583);
AND2_X1 g_g5585 (g4741, g4841, g5585);
AND2_X1 g_g5588 (g3028, g4969, g5588);
AND2_X1 g_g5593 (g4110, g4969, g5593);
AND2_X1 g_g5599 (g4745, g4969, g5599);
AND2_X1 g_g5624 (g5140, g2794, g5624);
AND2_X1 g_g5699 (g1667, g4841, g5699);
AND2_X1 g_g5700 (g1638, g4969, g5700);
AND2_X1 g_g5714 (g1532, g4733, g5714);
AND2_X1 g_g5765 (g1695, g5428, g5765);
AND2_X1 g_g5767 (g5344, g3079, g5767);
AND2_X1 g_g5783 (g1897, g5287, g5783);
AND2_X1 g_g5817 (g5395, g3091, g5817);
AND2_X1 g_g5894 (g1118, g5552, g5894);
AND2_X1 g_g5937 (g5562, g2407, g5937);
AND2_X1 g_g5969 (g5564, g2424, g5969);
AND2_X1 g_g5970 (g5605, g2424, g5970);
AND2_X1 g_g5984 (g1041, g5484, g5984);
AND2_X1 g_g6001 (g5540, g2407, g6001);
AND2_X1 g_g6002 (g5539, g2407, g6002);
AND3_X1 g_I10597 (g3769, g3754, g3735, I10597);
AND3_X1 g_g6003 (g3716, g5633, I10597, g6003);
AND2_X1 g_g6005 (g5557, g2407, g6005);
AND2_X1 g_g6006 (g5575, g2424, g6006);
AND2_X1 g_g6013 (g5589, g2424, g6013);
AND2_X1 g_g6021 (g5594, g2424, g6021);
AND2_X1 g_g6022 (g5595, g2424, g6022);
AND2_X1 g_g6039 (g1037, g5574, g6039);
AND2_X1 g_g6040 (g1462, g5578, g6040);
AND2_X1 g_g6041 (g5189, g4969, g6041);
AND2_X1 g_g6042 (g1041, g5581, g6042);
AND2_X1 g_g6043 (g1069, g5582, g6043);
AND2_X1 g_g6044 (g1467, g5584, g6044);
AND2_X1 g_g6045 (g1472, g5591, g6045);
AND2_X1 g_g6046 (g1073, g5592, g6046);
AND2_X1 g_g6047 (g1477, g5596, g6047);
AND2_X1 g_g6049 (g1045, g5597, g6049);
AND2_X1 g_g6052 (g1049, g5604, g6052);
AND2_X1 g_g6053 (g1053, g5608, g6053);
AND2_X1 g_g6054 (g1057, g5611, g6054);
AND2_X1 g_g6055 (g5239, g4202, g6055);
AND3_X1 g_g6056 (g3760, g5286, g1695, g6056);
AND2_X1 g_g6057 (g1061, g5617, g6057);
AND2_X1 g_g6058 (g5561, g3501, g6058);
AND2_X1 g_g6060 (g1065, g5623, g6060);
AND2_X1 g_g6061 (g5257, g1616, g6061);
AND2_X1 g_g6091 (g5712, g5038, g6091);
AND2_X1 g_g6098 (g5681, g1247, g6098);
AND2_X1 g_g6105 (g5618, g2817, g6105);
AND2_X1 g_g6107 (g5478, g1849, g6107);
AND2_X1 g_g6109 (g5453, g5335, g6109);
AND3_X1 g_g6112 (g5673, g4841, g5541, g6112);
AND2_X1 g_g6125 (g5548, g4202, g6125);
AND2_X1 g_g6145 (g1489, g5705, g6145);
AND2_X1 g_g6151 (g1494, g5709, g6151);
AND2_X1 g_g6154 (g1499, g5713, g6154);
AND2_X1 g_g6157 (g1130, g5717, g6157);
AND2_X1 g_g6160 (g1504, g5718, g6160);
AND2_X1 g_g6162 (g1134, g5724, g6162);
AND2_X1 g_g6166 (g1509, g5725, g6166);
AND2_X1 g_g6168 (g1138, g5191, g6168);
AND2_X1 g_g6171 (g5363, g4841, g6171);
AND2_X1 g_g6172 (g1514, g5192, g6172);
AND2_X1 g_g6175 (g4332, g5614, g6175);
AND2_X1 g_g6176 (g1149, g5198, g6176);
AND2_X1 g_g6182 (g1519, g5199, g6182);
AND2_X1 g_g6196 (g4927, g5615, g6196);
AND2_X1 g_g6204 (g5542, g5294, g6204);
AND2_X1 g_g6239 (g1514, g5314, g6239);
AND2_X1 g_g6266 (g1481, g5285, g6266);
AND2_X1 g_g6268 (g1092, g5309, g6268);
AND2_X1 g_g6394 (g5988, g5494, g6394);
AND2_X1 g_g6395 (g2157, g6007, g6395);
AND2_X1 g_g6396 (g661, g6008, g6396);
AND2_X1 g_g6399 (g5971, g5494, g6399);
AND2_X1 g_g6400 (g150, g6011, g6400);
AND2_X1 g_g6401 (g5971, g5367, g6401);
AND2_X1 g_g6402 (g665, g6012, g6402);
AND2_X1 g_g6405 (g5956, g5494, g6405);
AND2_X1 g_g6406 (g154, g6018, g6406);
AND2_X1 g_g6407 (g5956, g5367, g6407);
AND2_X1 g_g6408 (g669, g6019, g6408);
AND2_X1 g_g6409 (g706, g6020, g6409);
AND2_X1 g_g6411 (g5918, g5494, g6411);
AND2_X1 g_g6412 (g158, g6024, g6412);
AND2_X1 g_g6413 (g5939, g5367, g6413);
AND2_X1 g_g6414 (g673, g6025, g6414);
AND2_X1 g_g6415 (g5988, g5367, g6415);
AND2_X1 g_g6416 (g710, g6026, g6416);
AND2_X1 g_g6417 (g718, g6027, g6417);
AND2_X1 g_g6418 (g5897, g5494, g6418);
AND2_X1 g_g6419 (g162, g6032, g6419);
AND2_X1 g_g6420 (g5918, g5367, g6420);
AND2_X1 g_g6421 (g5847, g5384, g6421);
AND2_X1 g_g6422 (g714, g6033, g6422);
AND2_X1 g_g6423 (g5897, g5384, g6423);
AND2_X1 g_g6428 (g5874, g5494, g6428);
AND2_X1 g_g6429 (g168, g6035, g6429);
AND2_X1 g_g6430 (g5874, g5384, g6430);
AND2_X1 g_g6431 (g5847, g5494, g6431);
AND2_X1 g_g6433 (g778, g6134, g6433);
AND2_X1 g_g6434 (g855, g6048, g6434);
AND2_X1 g_g6437 (g859, g6050, g6437);
AND2_X1 g_g6438 (g4829, g6051, g6438);
AND2_X1 g_g6439 (g789, g6150, g6439);
AND2_X1 g_g6444 (g1676, g6125, g6444);
AND2_X1 g_g6447 (g734, g6073, g6447);
AND2_X1 g_g6448 (g5918, g5384, g6448);
AND2_X1 g_g6456 (g6116, g2407, g6456);
AND2_X1 g_g6460 (g6178, g2424, g6460);
AND2_X1 g_g6462 (g6215, g2424, g6462);
AND2_X1 g_g6464 (g6177, g2424, g6464);
AND2_X1 g_g6474 (g6203, g2424, g6474);
AND2_X1 g_g6487 (g5750, g4969, g6487);
AND2_X1 g_g6541 (g6144, g3510, g6541);
AND2_X1 g_g6554 (g5762, g1616, g6554);
AND2_X1 g_g6567 (g6265, g2424, g6567);
AND2_X1 g_g6574 (g1045, g5984, g6574);
AND2_X1 g_g6577 (g6142, g4160, g6577);
AND2_X1 g_g6578 (g6218, g3913, g6578);
AND2_X1 g_g6582 (g1122, g5894, g6582);
AND2_X1 g_g6611 (g3390, g6249, g6611);
AND2_X1 g_g6629 (g6023, g4841, g6629);
AND2_X1 g_g6633 (g5526, g5987, g6633);
AND2_X1 g_g6638 (g174, g5755, g6638);
AND2_X1 g_g6641 (g5939, g5494, g6641);
AND2_X1 g_g6643 (g1860, g5868, g6643);
AND2_X1 g_g6689 (g1519, g6239, g6689);
AND2_X1 g_g6715 (g677, g5843, g6715);
AND2_X1 g_g6726 (g5897, g5367, g6726);
AND2_X1 g_g6727 (g681, g5846, g6727);
AND2_X1 g_g6732 (g5874, g5367, g6732);
AND2_X1 g_g6733 (g685, g5873, g6733);
AND2_X1 g_g6738 (g5847, g5367, g6738);
AND2_X1 g_g6743 (g730, g5916, g6743);
AND2_X1 g_g6745 (g1872, g6198, g6745);
AND2_X1 g_g6753 (g5939, g5384, g6753);
AND2_X1 g_g6757 (g5874, g5412, g6757);
AND2_X1 g_g6762 (g5847, g5412, g6762);
AND2_X1 g_g6771 (g146, g6004, g6771);
AND2_X1 g_g6908 (g6478, g5246, g6908);
AND2_X1 g_g6914 (g6483, g5246, g6914);
AND2_X1 g_g6915 (g6493, g5246, g6915);
AND2_X1 g_g6916 (g727, g6515, g6916);
AND2_X1 g_g6923 (g6570, g5612, g6923);
AND2_X1 g_g6941 (g1126, g6582, g6941);
AND2_X1 g_g6949 (g5483, g6589, g6949);
AND2_X1 g_g6951 (g5511, g6595, g6951);
AND2_X1 g_g6954 (g5518, g6601, g6954);
AND2_X1 g_g6965 (g55, g6489, g6965);
AND2_X1 g_g6966 (g6580, g5580, g6966);
AND2_X1 g_g6970 (g5035, g6490, g6970);
AND2_X1 g_g6971 (g6424, g4969, g6971);
AND2_X1 g_g6972 (g5661, g6498, g6972);
AND2_X1 g_g6974 (g3613, g6505, g6974);
AND2_X1 g_g6976 (g4399, g6508, g6976);
AND2_X1 g_g6979 (g5095, g6511, g6979);
AND2_X1 g_g6990 (g799, g6517, g6990);
AND2_X1 g_g6991 (g5689, g6520, g6991);
AND2_X1 g_g6992 (g6610, g3519, g6992);
AND2_X1 g_g6994 (g3658, g6538, g6994);
AND2_X1 g_g6995 (g6435, g1616, g6995);
AND2_X1 g_g6996 (g3678, g6552, g6996);
AND2_X1 g_g6998 (g4474, g6555, g6998);
AND2_X1 g_g6999 (g815, g6556, g6999);
AND2_X1 g_g7001 (g3722, g6562, g7001);
AND2_X1 g_g7002 (g6770, g5054, g7002);
AND2_X1 g_g7003 (g1462, g6689, g7003);
AND2_X1 g_g7007 (g6627, g5072, g7007);
AND2_X1 g_g7008 (g6615, g5083, g7008);
AND2_X1 g_g7010 (g1049, g6574, g7010);
AND2_X1 g_g7017 (g3390, g6706, g7017);
AND2_X1 g_g7021 (g3390, g6673, g7021);
AND2_X1 g_g7027 (g3390, g6698, g7027);
AND2_X1 g_g7030 (g6705, g5723, g7030);
AND2_X1 g_g7031 (g3390, g6717, g7031);
AND2_X1 g_g7033 (g6716, g5190, g7033);
AND2_X1 g_g7036 (g6728, g5197, g7036);
AND2_X1 g_g7038 (g6466, g4841, g7038);
AND2_X1 g_g7041 (g6734, g5206, g7041);
AND2_X1 g_g7071 (g6639, g1872, g7071);
AND2_X1 g_g7079 (g4259, g6677, g7079);
AND2_X1 g_g7087 (g6440, g5311, g7087);
AND2_X1 g_g7096 (g6677, g5101, g7096);
AND2_X1 g_g7128 (g6926, g3047, g7128);
AND2_X1 g_g7136 (g4057, g6953, g7136);
AND2_X1 g_g7175 (g6893, g4841, g7175);
AND2_X1 g_g7177 (g7016, g5586, g7177);
AND2_X1 g_g7179 (g6121, g7035, g7179);
AND2_X1 g_g7181 (g6124, g7039, g7181);
AND2_X1 g_g7182 (g6902, g4969, g7182);
AND2_X1 g_g7183 (g6132, g7042, g7183);
AND2_X1 g_g7184 (g6138, g7043, g7184);
AND2_X1 g_g7186 (g6600, g7044, g7186);
AND2_X1 g_g7192 (g7026, g3526, g7192);
AND2_X1 g_g7193 (g6911, g1616, g7193);
AND2_X1 g_g7195 (g6984, g4226, g7195);
AND2_X1 g_g7197 (g7093, g5055, g7197);
AND2_X1 g_g7199 (g1467, g7003, g7199);
AND2_X1 g_g7212 (g1053, g7010, g7212);
AND2_X1 g_g7215 (g6111, g6984, g7215);
AND2_X1 g_g7217 (g1142, g6941, g7217);
AND2_X1 g_g7228 (g6688, g7090, g7228);
AND2_X1 g_g7232 (g6694, g7091, g7232);
AND2_X1 g_g7235 (g6699, g7094, g7235);
AND2_X1 g_g7238 (g6707, g7098, g7238);
AND2_X1 g_g7240 (g6719, g6894, g7240);
AND2_X1 g_g7242 (g7081, g6899, g7242);
AND2_X1 g_g7252 (g3591, g6977, g7252);
AND2_X1 g_g7271 (g6436, g6922, g7271);
AND2_X1 g_g7278 (g6965, g1745, g7278);
AND2_X1 g_g7282 (g5830, g6939, g7282);
AND2_X1 g_g7323 (g4065, g7171, g7323);
AND2_X1 g_g7412 (g7121, g4841, g7412);
AND2_X1 g_g7415 (g7222, g5603, g7415);
AND2_X1 g_g7416 (g7140, g4969, g7416);
AND2_X1 g_g7417 (g7144, g1616, g7417);
AND2_X1 g_g7419 (g7230, g3530, g7419);
AND2_X1 g_g7427 (g1472, g7199, g7427);
AND2_X1 g_g7429 (g1057, g7212, g7429);
AND2_X1 g_g7449 (g7272, g6901, g7449);
AND2_X1 g_g7536 (g4414, g7367, g7536);
AND2_X1 g_g7537 (g7363, g7411, g7537);
AND2_X1 g_g7552 (g7319, g5749, g7552);
AND2_X1 g_g7553 (g7367, g4135, g7553);
AND2_X1 g_g7554 (g7367, g4139, g7554);
AND2_X1 g_g7557 (g7367, g4147, g7557);
AND2_X1 g_g7559 (g7367, g4155, g7559);
AND2_X1 g_g7561 (g7367, g4163, g7561);
AND2_X1 g_g7564 (g7367, g4172, g7564);
AND2_X1 g_g7596 (g7428, g7028, g7596);
AND2_X1 g_g7597 (g7316, g4841, g7597);
AND2_X1 g_g7598 (g7483, g3466, g7598);
AND2_X1 g_g7600 (g7460, g3466, g7600);
AND2_X1 g_g7602 (g7476, g3466, g7602);
AND2_X1 g_g7604 (g7456, g3466, g7604);
AND2_X1 g_g7605 (g7435, g5607, g7605);
AND2_X1 g_g7606 (g7471, g3466, g7606);
AND2_X1 g_g7607 (g7325, g4969, g7607);
AND2_X1 g_g7608 (g7367, g4169, g7608);
AND2_X1 g_g7609 (g7467, g3466, g7609);
AND2_X1 g_g7611 (g7367, g4507, g7611);
AND2_X1 g_g7614 (g7367, g4176, g7614);
AND2_X1 g_g7615 (g7488, g3466, g7615);
AND2_X1 g_g7616 (g7367, g4517, g7616);
AND2_X1 g_g7625 (g7367, g4182, g7625);
AND2_X1 g_g7626 (g7463, g3466, g7626);
AND2_X1 g_g7628 (g7367, g4532, g7628);
AND2_X1 g_g7631 (g7367, g4187, g7631);
AND2_X1 g_g7632 (g7445, g3548, g7632);
AND2_X1 g_g7634 (g7367, g4549, g7634);
AND2_X1 g_g7652 (g7367, g4194, g7652);
AND2_X1 g_g7653 (g7480, g5754, g7653);
AND2_X1 g_g7654 (g7367, g4142, g7654);
AND2_X1 g_g7657 (g7367, g4201, g7657);
AND2_X1 g_g7658 (g7367, g4150, g7658);
AND2_X1 g_g7676 (g7367, g4216, g7676);
AND2_X1 g_g7677 (g7503, g5073, g7677);
AND2_X1 g_g7678 (g7367, g4158, g7678);
AND2_X1 g_g7679 (g7447, g5084, g7679);
AND2_X1 g_g7680 (g7367, g4166, g7680);
AND2_X1 g_g7681 (g7444, g5099, g7681);
AND2_X1 g_g7683 (g1061, g7429, g7683);
AND2_X1 g_g7689 (g7367, g4417, g7689);
AND2_X1 g_g7691 (g7367, g4427, g7691);
AND2_X1 g_g7692 (g7367, g4430, g7692);
AND2_X1 g_g7693 (g7367, g4445, g7693);
AND2_X1 g_g7694 (g7367, g4448, g7694);
AND2_X1 g_g7695 (g7367, g4466, g7695);
AND2_X1 g_g7696 (g7367, g4469, g7696);
AND2_X1 g_g7698 (g7367, g4483, g7698);
AND2_X1 g_g7699 (g7367, g4486, g7699);
AND2_X1 g_g7700 (g7367, g4494, g7700);
AND2_X1 g_g7701 (g7367, g4497, g7701);
AND2_X1 g_g7703 (g7367, g4504, g7703);
AND2_X1 g_g7705 (g7367, g4514, g7705);
AND2_X1 g_g7709 (g7367, g4529, g7709);
AND2_X1 g_g7713 (g4403, g7367, g7713);
AND2_X1 g_g7724 (g7337, g5938, g7724);
AND2_X1 g_g7827 (g7575, g7173, g7827);
AND2_X1 g_g7832 (g5343, g7599, g7832);
AND2_X1 g_g7833 (g6461, g7601, g7833);
AND2_X1 g_g7837 (g6470, g7610, g7837);
AND2_X1 g_g8059 (g7682, g7032, g8059);
AND2_X1 g_g8060 (g7535, g4841, g8060);
AND2_X1 g_g8062 (g7476, g7634, g8062);
AND2_X1 g_g8064 (g7483, g7634, g8064);
AND2_X1 g_g8066 (g7488, g7634, g8066);
AND2_X1 g_g8068 (g7687, g5610, g8068);
AND2_X1 g_g8069 (g7456, g7634, g8069);
AND2_X1 g_g8070 (g863, g7616, g8070);
AND2_X1 g_g8071 (g7540, g4969, g8071);
AND2_X1 g_g8074 (g855, g7616, g8074);
AND2_X1 g_g8075 (g7460, g7634, g8075);
AND2_X1 g_g8076 (g7690, g3521, g8076);
AND2_X1 g_g8077 (g859, g7616, g8077);
AND2_X1 g_g8078 (g7463, g7634, g8078);
AND2_X1 g_g8079 (g831, g7658, g8079);
AND2_X1 g_g8080 (g7467, g7634, g8080);
AND2_X1 g_g8081 (g834, g7658, g8081);
AND2_X1 g_g8087 (g7471, g7634, g8087);
AND2_X1 g_g8088 (g837, g7658, g8088);
AND2_X1 g_g8089 (g840, g7658, g8089);
AND2_X1 g_g8090 (g843, g7658, g8090);
AND2_X1 g_g8147 (g1065, g7683, g8147);
AND2_X1 g_g8150 (g846, g7658, g8150);
AND2_X1 g_g8151 (g849, g7658, g8151);
AND2_X1 g_g8153 (g852, g7658, g8153);
AND2_X1 g_g8229 (g8180, g5680, g8229);
AND2_X1 g_g8237 (g89, g8131, g8237);
AND2_X1 g_g8238 (g100, g8131, g8238);
AND2_X1 g_g8256 (g95, g8131, g8256);
AND2_X1 g_g8257 (g146, g8042, g8257);
AND2_X1 g_g8258 (g142, g8111, g8258);
AND2_X1 g_g8259 (g4538, g7855, g8259);
AND2_X1 g_g8260 (g138, g8111, g8260);
AND2_X1 g_g8261 (g174, g8042, g8261);
AND2_X1 g_g8262 (g4554, g7855, g8262);
AND2_X1 g_g8263 (g4555, g7905, g8263);
AND2_X1 g_g8264 (g105, g8131, g8264);
AND2_X1 g_g8265 (g134, g8111, g8265);
AND2_X1 g_g8266 (g2157, g8042, g8266);
AND2_X1 g_g8267 (g154, g8042, g8267);
AND2_X1 g_g8268 (g4568, g7905, g8268);
AND2_X1 g_g8269 (g4569, g7951, g8269);
AND2_X1 g_g8270 (g110, g8131, g8270);
AND2_X1 g_g8271 (g130, g8111, g8271);
AND2_X1 g_g8272 (g158, g8042, g8272);
AND2_X1 g_g8273 (g185, g8156, g8273);
AND2_X1 g_g8274 (g4580, g7951, g8274);
AND2_X1 g_g8275 (g4581, g7993, g8275);
AND2_X1 g_g8276 (g150, g8042, g8276);
AND2_X1 g_g8277 (g162, g8042, g8277);
AND2_X1 g_g8278 (g4589, g7993, g8278);
AND2_X1 g_g8280 (g114, g8111, g8280);
AND2_X1 g_g8281 (g168, g8042, g8281);
AND2_X1 g_g8282 (g179, g8156, g8282);
AND2_X1 g_g8283 (g267, g7838, g8283);
AND2_X1 g_g8285 (g118, g8111, g8285);
AND2_X1 g_g8286 (g180, g8156, g8286);
AND2_X1 g_g8287 (g4500, g7855, g8287);
AND2_X1 g_g8288 (g270, g7838, g8288);
AND2_X1 g_g8289 (g348, g7870, g8289);
AND2_X1 g_g8290 (g588, g8181, g8290);
AND2_X1 g_g8291 (g122, g8111, g8291);
AND2_X1 g_g8292 (g181, g8156, g8292);
AND2_X1 g_g8293 (g4510, g7855, g8293);
AND2_X1 g_g8294 (g281, g7838, g8294);
AND2_X1 g_g8295 (g4512, g7905, g8295);
AND2_X1 g_g8296 (g351, g7870, g8296);
AND2_X1 g_g8297 (g429, g7920, g8297);
AND2_X1 g_g8298 (g553, g8181, g8298);
AND2_X1 g_g8299 (g591, g8181, g8299);
AND2_X1 g_g8300 (g126, g8111, g8300);
AND2_X1 g_g8301 (g182, g8156, g8301);
AND2_X1 g_g8302 (g4521, g7855, g8302);
AND2_X1 g_g8303 (g284, g7838, g8303);
AND2_X1 g_g8304 (g4523, g7905, g8304);
AND2_X1 g_g8305 (g362, g7870, g8305);
AND2_X1 g_g8306 (g4525, g7951, g8306);
AND2_X1 g_g8307 (g432, g7920, g8307);
AND2_X1 g_g8308 (g510, g7966, g8308);
AND2_X1 g_g8309 (g550, g8181, g8309);
AND2_X1 g_g8310 (g573, g8181, g8310);
AND2_X1 g_g8311 (g4540, g7905, g8311);
AND2_X1 g_g8312 (g365, g7870, g8312);
AND2_X1 g_g8313 (g4542, g7951, g8313);
AND2_X1 g_g8314 (g443, g7920, g8314);
AND2_X1 g_g8315 (g4544, g7993, g8315);
AND2_X1 g_g8316 (g513, g7966, g8316);
AND2_X1 g_g8317 (g547, g8181, g8317);
AND2_X1 g_g8318 (g183, g8156, g8318);
AND2_X1 g_g8319 (g255, g7838, g8319);
AND2_X1 g_g8320 (g4557, g7951, g8320);
AND2_X1 g_g8321 (g446, g7920, g8321);
AND2_X1 g_g8322 (g4559, g7993, g8322);
AND2_X1 g_g8323 (g524, g7966, g8323);
AND2_X1 g_g8325 (g184, g8156, g8325);
AND2_X1 g_g8326 (g258, g7838, g8326);
AND2_X1 g_g8327 (g336, g7870, g8327);
AND2_X1 g_g8328 (g4571, g7993, g8328);
AND2_X1 g_g8329 (g527, g7966, g8329);
AND2_X1 g_g8330 (g261, g7838, g8330);
AND2_X1 g_g8331 (g339, g7870, g8331);
AND2_X1 g_g8332 (g417, g7920, g8332);
AND2_X1 g_g8333 (g563, g8181, g8333);
AND2_X1 g_g8334 (g264, g7838, g8334);
AND2_X1 g_g8335 (g342, g7870, g8335);
AND2_X1 g_g8336 (g420, g7920, g8336);
AND2_X1 g_g8337 (g498, g7966, g8337);
AND2_X1 g_g8338 (g570, g8181, g8338);
AND2_X1 g_g8339 (g345, g7870, g8339);
AND2_X1 g_g8340 (g423, g7920, g8340);
AND2_X1 g_g8341 (g501, g7966, g8341);
AND2_X1 g_g8359 (g642, g7793, g8359);
AND2_X1 g_g8361 (g426, g7920, g8361);
AND2_X1 g_g8362 (g504, g7966, g8362);
AND2_X1 g_g8377 (g507, g7966, g8377);
AND2_X1 g_g8378 (g677, g7887, g8378);
AND2_X1 g_g8379 (g691, g7793, g8379);
AND2_X1 g_g8380 (g681, g7887, g8380);
AND2_X1 g_g8382 (g685, g7887, g8382);
AND2_X1 g_g8383 (g730, g7937, g8383);
AND2_X1 g_g8384 (g636, g7793, g8384);
AND2_X1 g_g8385 (g695, g7811, g8385);
AND2_X1 g_g8403 (g639, g7793, g8403);
AND2_X1 g_g8404 (g710, g7937, g8404);
AND2_X1 g_g8405 (g741, g8018, g8405);
AND2_X1 g_g8438 (g649, g7793, g8438);
AND2_X1 g_g8439 (g699, g7811, g8439);
AND2_X1 g_g8440 (g714, g7937, g8440);
AND2_X1 g_g8441 (g746, g8018, g8441);
AND2_X1 g_g8455 (g652, g7793, g8455);
AND2_X1 g_g8456 (g703, g7811, g8456);
AND2_X1 g_g8457 (g724, g7811, g8457);
AND2_X1 g_g8458 (g756, g8199, g8458);
AND2_X1 g_g8459 (g655, g7793, g8459);
AND2_X1 g_g8460 (g757, g8199, g8460);
AND2_X1 g_g8461 (g658, g7793, g8461);
AND2_X1 g_g8462 (g49, g8199, g8462);
AND2_X1 g_g8513 (g718, g7937, g8513);
AND2_X1 g_g8542 (g661, g7887, g8542);
AND2_X1 g_g8543 (g706, g7887, g8543);
AND2_X1 g_g8584 (g8146, g7034, g8584);
AND2_X1 g_g8607 (g8154, g5616, g8607);
AND2_X1 g_g8609 (g7828, g4969, g8609);
AND2_X1 g_g8610 (g665, g7887, g8610);
AND2_X1 g_g8611 (g669, g7887, g8611);
AND2_X1 g_g8612 (g673, g7887, g8612);
AND2_X1 g_g8620 (g751, g8199, g8620);
AND2_X1 g_g8621 (g734, g7937, g8621);
AND2_X1 g_g8622 (g738, g7811, g8622);
AND2_X1 g_g8623 (g755, g8199, g8623);
AND2_X1 g_g8624 (g754, g8199, g8624);
AND2_X1 g_g8626 (g752, g8199, g8626);
AND2_X1 g_g8628 (g753, g8199, g8628);
AND2_X1 g_g8643 (g547, g8094, g8643);
AND2_X1 g_g8645 (g550, g8094, g8645);
AND2_X1 g_g8646 (g553, g8094, g8646);
AND2_X1 g_g8648 (g588, g8094, g8648);
AND2_X1 g_g8650 (g591, g8094, g8650);
AND2_X1 g_g8652 (g563, g8094, g8652);
AND2_X1 g_g8653 (g573, g8094, g8653);
AND2_X1 g_g8654 (g570, g8094, g8654);
AND2_X1 g_g8660 (g1069, g8147, g8660);
AND2_X1 g_g8686 (g3819, g8342, g8686);
AND2_X1 g_g8687 (g3488, g8363, g8687);
AND2_X1 g_g8688 (g3812, g8342, g8688);
AND2_X1 g_g8690 (g3485, g8363, g8690);
AND2_X1 g_g8691 (g3805, g8342, g8691);
AND2_X1 g_g8692 (g3462, g8363, g8692);
AND2_X1 g_g8693 (g3798, g8342, g8693);
AND2_X1 g_g8695 (g2709, g8363, g8695);
AND2_X1 g_g8696 (g3743, g8342, g8696);
AND2_X1 g_g8697 (g3761, g8342, g8697);
AND2_X1 g_g8698 (g3774, g8342, g8698);
AND2_X1 g_g8700 (g3784, g8342, g8700);
AND2_X1 g_g8701 (g2700, g8363, g8701);
AND2_X1 g_g8702 (g2837, g8386, g8702);
AND2_X1 g_g8703 (g3574, g8407, g8703);
AND2_X1 g_g8704 (g2829, g8386, g8704);
AND2_X1 g_g8705 (g2798, g8421, g8705);
AND2_X1 g_g8708 (g3557, g8407, g8708);
AND2_X1 g_g8709 (g2818, g8386, g8709);
AND2_X1 g_g8710 (g2790, g8421, g8710);
AND2_X1 g_g8711 (g3542, g8407, g8711);
AND2_X1 g_g8712 (g2804, g8386, g8712);
AND2_X1 g_g8713 (g2777, g8421, g8713);
AND2_X1 g_g8714 (g2873, g8407, g8714);
AND2_X1 g_g8715 (g2761, g8386, g8715);
AND2_X1 g_g8716 (g3506, g8443, g8716);
AND2_X1 g_g8717 (g2764, g8421, g8717);
AND2_X1 g_g8718 (g2774, g8386, g8718);
AND2_X1 g_g8719 (g2821, g8443, g8719);
AND2_X1 g_g8720 (g3825, g8421, g8720);
AND2_X1 g_g8721 (g2703, g8464, g8721);
AND2_X1 g_g8722 (g2787, g8386, g8722);
AND2_X1 g_g8723 (g2706, g8421, g8723);
AND2_X1 g_g8724 (g3822, g8464, g8724);
AND2_X1 g_g8725 (g3008, g8493, g8725);
AND2_X1 g_g8726 (g2795, g8386, g8726);
AND2_X1 g_g8727 (g2724, g8421, g8727);
AND2_X1 g_g8728 (g3815, g8464, g8728);
AND2_X1 g_g8729 (g2999, g8493, g8729);
AND2_X1 g_g8730 (g2863, g8407, g8730);
AND2_X1 g_g8731 (g2743, g8421, g8731);
AND2_X1 g_g8732 (g3808, g8464, g8732);
AND2_X1 g_g8733 (g2996, g8493, g8733);
AND2_X1 g_g8735 (g2807, g8443, g8735);
AND2_X1 g_g8736 (g3771, g8464, g8736);
AND2_X1 g_g8737 (g2992, g8493, g8737);
AND2_X1 g_g8738 (g8619, g3338, g8738);
AND2_X1 g_g8739 (g3780, g8464, g8739);
AND2_X1 g_g8740 (g2966, g8493, g8740);
AND2_X1 g_g8741 (g3787, g8464, g8741);
AND2_X1 g_g8742 (g2973, g8493, g8742);
AND2_X1 g_g8744 (g3802, g8464, g8744);
AND2_X1 g_g8745 (g2982, g8493, g8745);
AND2_X1 g_g8748 (g2721, g8483, g8748);
AND2_X1 g_g8749 (g2989, g8493, g8749);
AND2_X1 g_g8764 (g8231, g4969, g8764);
AND2_X1 g_g8779 (g8634, g7037, g8779);
AND2_X1 g_g8793 (g8637, g5622, g8793);
AND2_X1 g_g8813 (g255, g8524, g8813);
AND2_X1 g_g8814 (g3880, g8463, g8814);
AND2_X1 g_g8815 (g258, g8524, g8815);
AND2_X1 g_g8816 (g336, g8545, g8816);
AND2_X1 g_g8817 (g4545, g8482, g8817);
AND2_X1 g_g8820 (g261, g8524, g8820);
AND2_X1 g_g8821 (g339, g8545, g8821);
AND2_X1 g_g8822 (g417, g8564, g8822);
AND2_X1 g_g8823 (g4561, g8512, g8823);
AND2_X1 g_g8824 (g264, g8524, g8824);
AND2_X1 g_g8825 (g342, g8545, g8825);
AND2_X1 g_g8826 (g420, g8564, g8826);
AND2_X1 g_g8827 (g498, g8585, g8827);
AND2_X1 g_g8828 (g4573, g8541, g8828);
AND2_X1 g_g8829 (g267, g8524, g8829);
AND2_X1 g_g8830 (g345, g8545, g8830);
AND2_X1 g_g8831 (g423, g8564, g8831);
AND2_X1 g_g8832 (g501, g8585, g8832);
AND2_X1 g_g8833 (g4583, g8562, g8833);
AND2_X1 g_g8835 (g270, g8524, g8835);
AND2_X1 g_g8836 (g348, g8545, g8836);
AND2_X1 g_g8837 (g426, g8564, g8837);
AND2_X1 g_g8838 (g504, g8585, g8838);
AND2_X1 g_g8839 (g4050, g8581, g8839);
AND2_X1 g_g8840 (g4590, g8582, g8840);
AND2_X1 g_g8841 (g351, g8545, g8841);
AND2_X1 g_g8842 (g429, g8564, g8842);
AND2_X1 g_g8843 (g507, g8585, g8843);
AND2_X1 g_g8844 (g4056, g8602, g8844);
AND2_X1 g_g8845 (g432, g8564, g8845);
AND2_X1 g_g8846 (g510, g8585, g8846);
AND2_X1 g_g8848 (g281, g8524, g8848);
AND2_X1 g_g8849 (g513, g8585, g8849);
AND2_X1 g_g8851 (g284, g8524, g8851);
AND2_X1 g_g8852 (g362, g8545, g8852);
AND2_X1 g_g8853 (g365, g8545, g8853);
AND2_X1 g_g8854 (g443, g8564, g8854);
AND2_X1 g_g8857 (g446, g8564, g8857);
AND2_X1 g_g8858 (g524, g8585, g8858);
AND2_X1 g_g8860 (g527, g8585, g8860);
AND2_X1 g_g8876 (g8769, g6102, g8876);
AND2_X1 g_g8877 (g8773, g6104, g8877);
AND2_X1 g_g8878 (g8777, g6106, g8878);
AND2_X1 g_g8879 (g8782, g6108, g8879);
AND2_X1 g_g8892 (g8681, g4969, g8892);
AND2_X1 g_g8901 (g8804, g5631, g8901);
AND2_X1 g_g8911 (g8798, g7688, g8911);
AND2_X1 g_g8912 (g8796, g8239, g8912);
AND2_X1 g_g8914 (g8795, g8239, g8914);
AND2_X1 g_g8915 (g8794, g8239, g8915);
AND2_X1 g_g8919 (g4567, g8743, g8919);
AND2_X1 g_g8920 (g4578, g8746, g8920);
AND2_X1 g_g8921 (g4579, g8747, g8921);
AND2_X1 g_g8922 (g4586, g8750, g8922);
AND2_X1 g_g8923 (g4587, g8751, g8923);
AND2_X1 g_g8924 (g4588, g8752, g8924);
AND2_X1 g_g8925 (g4592, g8754, g8925);
AND2_X1 g_g8926 (g4593, g8755, g8926);
AND2_X1 g_g8927 (g4594, g8756, g8927);
AND2_X1 g_g8928 (g4595, g8757, g8928);
AND2_X1 g_g8929 (g3865, g8759, g8929);
AND2_X1 g_g8930 (g3866, g8760, g8930);
AND2_X1 g_g8931 (g3867, g8761, g8931);
AND2_X1 g_g8932 (g3868, g8762, g8932);
AND2_X1 g_g8933 (g4511, g8765, g8933);
AND2_X1 g_g8934 (g3873, g8766, g8934);
AND2_X1 g_g8935 (g3874, g8767, g8935);
AND2_X1 g_g8936 (g3875, g8768, g8936);
AND2_X1 g_g8937 (g4524, g8770, g8937);
AND2_X1 g_g8938 (g3878, g8771, g8938);
AND2_X1 g_g8939 (g3879, g8772, g8939);
AND2_X1 g_g8940 (g4543, g8775, g8940);
AND2_X1 g_g8941 (g3882, g8776, g8941);
AND2_X1 g_g8942 (g4522, g8780, g8942);
AND2_X1 g_g8943 (g4560, g8781, g8943);
AND2_X1 g_g8944 (g4539, g8783, g8944);
AND2_X1 g_g8945 (g4541, g8784, g8945);
AND2_X1 g_g8946 (g4556, g8786, g8946);
AND2_X1 g_g8947 (g4558, g8787, g8947);
AND2_X1 g_g8948 (g4570, g8789, g8948);
AND2_X1 g_g8949 (g4572, g8790, g8949);
AND2_X1 g_g8950 (g4582, g8791, g8950);
AND2_X1 g_g8951 (g8785, g6072, g8951);
AND2_X1 g_g8952 (g8788, g6075, g8952);
AND2_X1 g_g8953 (g8758, g6093, g8953);
AND2_X1 g_g8954 (g8763, g6097, g8954);
AND2_X1 g_g8961 (g8885, g5317, g8961);
AND2_X1 g_g8962 (g8890, g5317, g8962);
AND2_X1 g_g8963 (g8891, g5317, g8963);
AND2_X1 g_g8976 (g8903, g6588, g8976);
AND2_X1 g_g8978 (g8909, g5587, g8978);
AND2_X1 g_g9012 (g8908, g8239, g9012);
AND2_X1 g_g9013 (g8907, g8239, g9013);
AND2_X1 g_g9014 (g8906, g8239, g9014);
AND2_X1 g_g9015 (g8905, g8239, g9015);
AND2_X1 g_g9016 (g8904, g8239, g9016);
AND2_X1 g_g9021 (g8886, g5317, g9021);
AND2_X1 g_g9022 (g8887, g5317, g9022);
AND2_X1 g_g9023 (g8888, g5317, g9023);
AND2_X1 g_g9024 (g8884, g5317, g9024);
AND2_X1 g_g9025 (g8889, g5317, g9025);
AND2_X1 g_g9037 (g8965, g5345, g9037);
AND2_X1 g_g9038 (g8966, g5345, g9038);
AND2_X1 g_g9080 (g9011, g5598, g9080);
AND2_X1 g_g9084 (g8964, g5345, g9084);
AND2_X1 g_g9118 (g9046, g5345, g9118);
AND2_X1 g_g9119 (g9049, g5345, g9119);
AND2_X1 g_g9120 (g9052, g5345, g9120);
AND2_X1 g_g9130 (g9054, g5345, g9130);
AND2_X1 g_g9131 (g9055, g5345, g9131);
AND2_X1 g_g9142 (g9124, g6059, g9142);
AND2_X1 g_g9143 (g9122, g6089, g9143);
AND2_X1 g_g9144 (g9123, g6096, g9144);
AND2_X1 g_g9146 (g9135, g6101, g9146);
AND2_X1 g_g9147 (g9136, g6103, g9147);
AND2_X1 g_g9158 (g9137, g6070, g9158);
AND2_X1 g_g9159 (g9138, g6074, g9159);
AND2_X1 g_g9160 (g9139, g6092, g9160);
AND2_X1 g_g9226 (g9220, g5403, g9226);
AND2_X1 g_g9238 (g4748, g9223, g9238);
AND2_X1 g_g9240 (g9223, g5261, g9240);
AND2_X1 g_g9247 (g4748, g9227, g9247);
AND2_X1 g_g9251 (g4748, g9230, g9251);
AND2_X1 g_g9258 (g9227, g5628, g9258);
AND2_X1 g_g9259 (g9230, g5639, g9259);
AND2_X1 g_g9270 (g4748, g9241, g9270);
AND2_X1 g_g9271 (g4748, g9244, g9271);
AND2_X1 g_g9272 (g4748, g9248, g9272);
AND2_X1 g_g9273 (g4748, g9252, g9273);
AND2_X1 g_g9274 (g4748, g9255, g9274);
AND2_X1 g_g9275 (g9241, g5645, g9275);
AND2_X1 g_g9276 (g9244, g5649, g9276);
AND2_X1 g_g9277 (g9248, g5654, g9277);
AND2_X1 g_g9278 (g9252, g5658, g9278);
AND2_X1 g_g9279 (g9255, g5665, g9279);
AND2_X1 g_g9327 (g9316, g5757, g9327);
AND2_X1 g_g9328 (g9324, g6465, g9328);
AND2_X1 g_g9334 (g9318, g6205, g9334);
AND2_X1 g_g9335 (g9320, g6206, g9335);
AND2_X1 g_g9343 (g9328, g1738, g9343);
AND2_X1 g_g9344 (g9329, g6211, g9344);
AND2_X1 g_g9345 (g9330, g6217, g9345);
AND2_X1 g_g9346 (g9331, g6222, g9346);
AND2_X1 g_g9347 (g9332, g6226, g9347);
AND2_X1 g_g9348 (g9333, g6229, g9348);
AND2_X1 g_g9349 (g9340, g5690, g9349);
AND2_X1 g_g9359 (g4748, g9340, g9359);
AND2_X1 g_g9371 (g9352, g5917, g9371);
AND2_X1 g_g9384 (g9383, g6245, g9384);
OR3_X1 g_g1690 (g1021, g1025, g1018, g1690);
OR4_X1 g_I5757 (g969, g970, g966, g963, I5757);
OR4_X1 g_g1872 (g971, g962, g972, I5757, g1872);
OR2_X1 g_g1955 (g1189, g16, g1955);
OR2_X1 g_g2043 (g1263, g1257, g2043);
OR4_X1 g_g2206 (g1363, g1364, g1365, g1366, g2206);
OR4_X1 g_g2213 (g1367, g1368, g1369, g1370, g2213);
OR4_X1 g_g2214 (g1376, g1377, g1378, g1379, g2214);
OR4_X1 g_g2229 (g1371, g1372, g1373, g1374, g2229);
OR4_X1 g_g2230 (g1380, g1381, g1382, g1383, g2230);
OR4_X1 g_g2262 (g1384, g1385, g1386, g1387, g2262);
OR4_X1 g_I6208 (g891, g896, g901, g906, I6208);
OR4_X1 g_I6209 (g911, g916, g921, g883, I6209);
OR2_X1 g_g2368 (I6208, I6209, g2368);
OR2_X1 g_g2845 (g1877, g576, g2845);
OR2_X1 g_g3097 (g1746, g287, g3097);
OR2_X1 g_g3131 (g1749, g368, g3131);
OR2_X1 g_g3160 (g1751, g449, g3160);
OR2_X1 g_g3192 (g1756, g530, g3192);
OR2_X1 g_g3339 (g1424, g2014, g3339);
OR2_X1 g_g3541 (g1663, g1421, g3541);
OR4_X1 g_I7232 (g2367, g2352, g2378, g2330, I7232);
OR4_X1 g_I7233 (g2315, g2385, g2294, g2395, I7233);
OR2_X1 g_g3760 (I7232, I7233, g3760);
OR2_X1 g_g3986 (g202, g3129, g3986);
OR2_X1 g_g4055 (g187, g3012, g4055);
OR2_X1 g_g4072 (g196, g2995, g4072);
OR2_X1 g_g4179 (g207, g3083, g4179);
OR2_X1 g_g4249 (g3617, g1639, g4249);
OR2_X1 g_g4264 (g2490, g3315, g4264);
OR4_X1 g_I8224 (g3019, g3029, g3038, g3052, I8224);
OR4_X1 g_I8225 (g3062, g2712, g2734, g2752, I8225);
OR2_X1 g_g4280 (I8224, I8225, g4280);
OR2_X1 g_g4283 (g3587, g2665, g4283);
OR2_X1 g_g4295 (g2828, g2668, g4295);
OR2_X1 g_g4297 (g3617, g3602, g4297);
OR2_X1 g_g4364 (g2952, g1725, g4364);
OR3_X1 g_I8363 (g2655, g1163, g1160, I8363);
OR4_X1 g_g4374 (g1182, g1186, g1179, I8363, g4374);
OR2_X1 g_g4413 (g2371, g3285, g4413);
OR2_X1 g_g4688 (g4193, g3190, g4688);
OR3_X1 g_I9029 (g4504, g4494, g4430, I9029);
OR4_X1 g_g4727 (g4417, g4172, g4163, I9029, g4727);
OR3_X1 g_I9038 (g4507, g4497, g4486, I9038);
OR3_X1 g_g4734 (g4469, g4448, I9038, g4734);
OR3_X1 g_I9041 (g4483, g4466, g4445, I9041);
OR4_X1 g_g4735 (g4427, g4414, g4403, I9041, g4735);
OR3_X1 g_I9044 (g4150, g4142, g4549, I9044);
OR3_X1 g_g4736 (g4532, g4517, I9044, g4736);
OR3_X1 g_I9047 (g4155, g4147, g4139, I9047);
OR4_X1 g_g4737 (g4135, g4529, g4514, I9047, g4737);
OR2_X1 g_g4747 (g3984, g2912, g4747);
OR3_X1 g_I9099 (g4127, g4123, g4117, I9099);
OR4_X1 g_g4786 (g4107, g4097, g4124, I9099, g4786);
OR4_X1 g_I9107 (g4133, g4145, g4138, g4132, I9107);
OR4_X1 g_g4790 (g4185, g4131, g4129, I9107, g4790);
OR2_X1 g_g4812 (g2490, g4237, g4812);
OR2_X1 g_g4829 (g863, g4051, g4829);
OR2_X1 g_g4870 (g4154, g3081, g4870);
OR2_X1 g_g4876 (g4159, g4167, g4876);
OR2_X1 g_g4927 (g4318, g1590, g4927);
OR2_X1 g_g5021 (g943, g4501, g5021);
OR2_X1 g_g5036 (g4047, g2972, g5036);
OR4_X1 g_g5040 (g3900, g3895, g3890, g4363, g5040);
OR2_X1 g_g5052 (g4049, g4054, g5052);
OR4_X1 g_g5057 (g3939, g3925, g3915, g3907, g5057);
OR2_X1 g_g5070 (g4052, g4058, g5070);
OR2_X1 g_g5138 (g4108, g3049, g5138);
OR2_X1 g_g5140 (g4333, g3509, g5140);
OR2_X1 g_g5188 (g5008, g4365, g5188);
OR2_X1 g_g5193 (g5017, g4366, g5193);
OR2_X1 g_g5194 (g5018, g4367, g5194);
OR2_X1 g_g5195 (g5019, g4368, g5195);
OR2_X1 g_g5196 (g5020, g4369, g5196);
OR2_X1 g_g5200 (g5029, g4375, g5200);
OR2_X1 g_g5201 (g5030, g4376, g5201);
OR2_X1 g_g5202 (g5031, g4377, g5202);
OR2_X1 g_g5203 (g5032, g4378, g5203);
OR2_X1 g_g5204 (g5033, g4379, g5204);
OR2_X1 g_g5205 (g5034, g4380, g5205);
OR2_X1 g_g5208 (g5043, g4383, g5208);
OR2_X1 g_g5209 (g5044, g4384, g5209);
OR2_X1 g_g5210 (g5045, g4385, g5210);
OR2_X1 g_g5211 (g5046, g4386, g5211);
OR2_X1 g_g5212 (g5047, g4387, g5212);
OR2_X1 g_g5213 (g5048, g4388, g5213);
OR2_X1 g_g5214 (g5049, g4389, g5214);
OR2_X1 g_g5215 (g5050, g4390, g5215);
OR2_X1 g_g5216 (g5062, g4391, g5216);
OR2_X1 g_g5217 (g5063, g4392, g5217);
OR2_X1 g_g5218 (g5064, g4393, g5218);
OR2_X1 g_g5219 (g5065, g4394, g5219);
OR2_X1 g_g5220 (g5066, g4395, g5220);
OR2_X1 g_g5221 (g5067, g4396, g5221);
OR2_X1 g_g5222 (g5068, g4397, g5222);
OR2_X1 g_g5223 (g5069, g4398, g5223);
OR2_X1 g_g5227 (g5077, g4407, g5227);
OR2_X1 g_g5228 (g5078, g4408, g5228);
OR2_X1 g_g5229 (g5079, g4409, g5229);
OR2_X1 g_g5230 (g5080, g4410, g5230);
OR2_X1 g_g5231 (g5081, g4411, g5231);
OR2_X1 g_g5232 (g5082, g4412, g5232);
OR2_X1 g_g5233 (g5089, g4420, g5233);
OR2_X1 g_g5234 (g5090, g4421, g5234);
OR2_X1 g_g5235 (g5091, g4422, g5235);
OR2_X1 g_g5236 (g5092, g4423, g5236);
OR2_X1 g_g5237 (g5093, g4424, g5237);
OR2_X1 g_g5238 (g5094, g4425, g5238);
OR2_X1 g_g5241 (g5104, g4433, g5241);
OR2_X1 g_g5242 (g5105, g4434, g5242);
OR2_X1 g_g5243 (g5106, g4435, g5243);
OR2_X1 g_g5244 (g5107, g4436, g5244);
OR2_X1 g_g5245 (g5108, g4437, g5245);
OR2_X1 g_g5253 (g5116, g4451, g5253);
OR2_X1 g_g5254 (g5117, g4452, g5254);
OR2_X1 g_g5255 (g5118, g4453, g5255);
OR2_X1 g_g5256 (g5119, g4454, g5256);
OR2_X1 g_g5259 (g5122, g4472, g5259);
OR2_X1 g_g5260 (g5123, g4473, g5260);
OR2_X1 g_g5264 (g5125, g4490, g5264);
OR2_X1 g_g5265 (g5126, g4491, g5265);
OR3_X1 g_g5317 (g4727, g4737, g4735, g5317);
OR2_X1 g_g5343 (g4690, g2862, g5343);
OR2_X1 g_g5345 (g4736, g4734, g5345);
OR2_X1 g_g5440 (g4790, g4786, g5440);
OR2_X1 g_g5483 (g4740, g4098, g5483);
OR2_X1 g_g5511 (g4743, g4109, g5511);
OR2_X1 g_g5518 (g4744, g4118, g5518);
OR2_X1 g_g5537 (g3617, g4835, g5537);
OR2_X1 g_g5545 (g3617, g4824, g5545);
OR2_X1 g_g5549 (g2935, g4712, g5549);
OR2_X1 g_g5561 (g4168, g4797, g5561);
OR2_X1 g_g5566 (g3617, g4810, g5566);
OR2_X1 g_g5572 (g5051, g1236, g5572);
OR2_X1 g_g5673 (g4823, g4872, g5673);
OR2_X1 g_g5698 (g5057, g5040, g5698);
OR2_X1 g_g5704 (g4936, g4334, g5704);
OR2_X1 g_g5706 (g4955, g4342, g5706);
OR2_X1 g_g5707 (g4956, g4343, g5707);
OR2_X1 g_g5708 (g2889, g4699, g5708);
OR2_X1 g_g5710 (g4958, g4351, g5710);
OR2_X1 g_g5711 (g4959, g4352, g5711);
OR2_X1 g_g5715 (g4961, g4355, g5715);
OR2_X1 g_g5716 (g4962, g4356, g5716);
OR2_X1 g_g5722 (g5001, g4361, g5722);
OR2_X1 g_g5830 (g5714, g5142, g5830);
OR2_X1 g_g6115 (g3617, g5558, g6115);
OR2_X1 g_g6116 (g5546, g4681, g6116);
OR2_X1 g_g6120 (g3617, g5555, g6120);
OR2_X1 g_g6121 (g5425, g4785, g6121);
OR2_X1 g_g6123 (g3617, g5556, g6123);
OR2_X1 g_g6124 (g5432, g4789, g6124);
OR2_X1 g_g6132 (g5436, g4793, g6132);
OR2_X1 g_g6138 (g5438, g5442, g6138);
OR2_X1 g_g6144 (g4175, g5458, g6144);
OR2_X1 g_g6249 (g4066, g5313, g6249);
OR2_X1 g_g6262 (g4074, g5334, g6262);
OR3_X1 g_g6270 (g1000, g5335, g1909, g6270);
OR2_X1 g_g6436 (g6266, g5699, g6436);
OR2_X1 g_g6440 (g6268, g5700, g6440);
OR2_X1 g_g6445 (g6105, g6107, g6445);
OR3_X1 g_g6457 (g6196, g6209, g4937, g6457);
OR4_X1 g_g6458 (g6184, g6259, g6174, g6214, g6458);
OR3_X1 g_I11603 (g6193, g6197, g6175, I11603);
OR3_X1 g_g6459 (g6259, g6185, I11603, g6459);
OR2_X1 g_g6470 (g5817, g2934, g6470);
OR2_X1 g_g6525 (g6112, g5547, g6525);
OR2_X1 g_g6543 (g6125, g1553, g6543);
OR3_X1 g_g6565 (g2396, g6131, g1603, g6565);
OR2_X1 g_g6579 (g6098, g1975, g6579);
OR2_X1 g_g6580 (g6039, g6041, g6580);
OR2_X1 g_g6585 (g3617, g6119, g6585);
OR2_X1 g_g6590 (g3617, g6153, g6590);
OR2_X1 g_g6600 (g5443, g6055, g6600);
OR2_X1 g_g6602 (g6058, g3092, g6602);
OR2_X1 g_g6610 (g4180, g6061, g6610);
OR2_X1 g_g6673 (g4053, g5937, g6673);
OR2_X1 g_g6685 (g4067, g5969, g6685);
OR2_X1 g_g6686 (g4068, g5970, g6686);
OR2_X1 g_g6688 (g6145, g5570, g6688);
OR2_X1 g_g6694 (g6151, g5573, g6694);
OR2_X1 g_g6698 (g4073, g6001, g6698);
OR2_X1 g_g6699 (g6154, g5579, g6699);
OR2_X1 g_g6705 (g6157, g5583, g6705);
OR2_X1 g_g6706 (g4077, g6002, g6706);
OR2_X1 g_g6707 (g6160, g5585, g6707);
OR2_X1 g_g6710 (g55, g6264, g6710);
OR2_X1 g_g6716 (g6162, g5588, g6716);
OR2_X1 g_g6717 (g4082, g6005, g6717);
OR2_X1 g_g6718 (g4083, g6006, g6718);
OR2_X1 g_g6719 (g6166, g6171, g6719);
OR2_X1 g_g6728 (g6168, g5593, g6728);
OR2_X1 g_g6734 (g6176, g5599, g6734);
OR2_X1 g_g6735 (g4091, g6013, g6735);
OR2_X1 g_g6739 (g4099, g6021, g6739);
OR2_X1 g_g6740 (g4100, g6022, g6740);
OR2_X1 g_g6906 (g6715, g6726, g6906);
OR2_X1 g_g6907 (g6727, g6732, g6907);
OR2_X1 g_g6912 (g4199, g6567, g6912);
OR2_X1 g_g6913 (g6733, g6738, g6913);
OR2_X1 g_g6917 (g6743, g6753, g6917);
OR2_X1 g_g6919 (g6771, g6394, g6919);
OR2_X1 g_g6920 (g6395, g6399, g6920);
OR2_X1 g_g6921 (g6396, g6401, g6921);
OR2_X1 g_g6924 (g6400, g6405, g6924);
OR2_X1 g_g6925 (g6402, g6407, g6925);
OR2_X1 g_g6926 (g6406, g6411, g6926);
OR2_X1 g_g6927 (g6408, g6413, g6927);
OR2_X1 g_g6928 (g6409, g6415, g6928);
OR2_X1 g_g6929 (g6412, g6418, g6929);
OR2_X1 g_g6930 (g6414, g6420, g6930);
OR2_X1 g_g6931 (g6416, g6421, g6931);
OR2_X1 g_g6932 (g6417, g6423, g6932);
OR2_X1 g_g6933 (g6419, g6428, g6933);
OR2_X1 g_g6934 (g6422, g6430, g6934);
OR2_X1 g_g6935 (g6429, g6431, g6935);
OR2_X1 g_g6952 (g6633, g6204, g6952);
OR2_X1 g_g6964 (g6447, g6448, g6964);
OR2_X1 g_g6980 (g6745, g6028, g6980);
OR2_X1 g_g7016 (g6042, g6487, g7016);
OR2_X1 g_g7020 (g3617, g6578, g7020);
OR2_X1 g_g7025 (g6541, g3095, g7025);
OR2_X1 g_g7026 (g4186, g6554, g7026);
OR2_X1 g_g7029 (g6433, g5765, g7029);
OR2_X1 g_g7040 (g6439, g5783, g7040);
OR2_X1 g_g7062 (g4048, g6456, g7062);
OR2_X1 g_g7080 (g4086, g6462, g7080);
OR2_X1 g_g7081 (g6172, g6629, g7081);
OR3_X1 g_g7083 (g5448, g6267, g6710, g7083);
OR2_X1 g_g7086 (g4101, g6464, g7086);
OR2_X1 g_g7088 (g6638, g6641, g7088);
OR2_X1 g_g7089 (g4128, g6474, g7089);
OR2_X1 g_g7165 (g6434, g6908, g7165);
OR2_X1 g_g7166 (g6437, g6914, g7166);
OR2_X1 g_g7167 (g6438, g6915, g7167);
OR2_X1 g_g7170 (g6916, g6444, g7170);
OR2_X1 g_g7191 (g7071, g6980, g7191);
OR2_X1 g_g7202 (g6028, g7071, g7202);
OR2_X1 g_g7220 (g1304, g7062, g7220);
OR2_X1 g_g7222 (g6049, g6971, g7222);
OR2_X1 g_g7227 (g6992, g3128, g7227);
OR2_X1 g_g7230 (g4190, g6995, g7230);
OR2_X1 g_g7248 (g7079, g5652, g7248);
OR2_X1 g_g7254 (g6923, g5298, g7254);
OR3_X1 g_I13220 (g58, g6258, g5418, I13220);
OR3_X1 g_g7258 (g7083, g5403, I13220, g7258);
OR2_X1 g_g7272 (g6182, g7038, g7272);
OR2_X1 g_g7337 (g7278, g4546, g7337);
OR2_X1 g_g7363 (g7136, g6903, g7363);
OR2_X1 g_g7421 (g6745, g7202, g7421);
OR3_X1 g_I13553 (g1166, g1167, g1170, I13553);
OR3_X1 g_g7426 (g1173, g7217, I13553, g7426);
OR2_X1 g_g7428 (g6040, g7175, g7428);
OR2_X1 g_g7435 (g6052, g7182, g7435);
OR2_X1 g_g7436 (g7183, g6975, g7436);
OR2_X1 g_g7438 (g7184, g6978, g7438);
OR2_X1 g_g7443 (g7192, g3158, g7443);
OR2_X1 g_g7445 (g4192, g7193, g7445);
OR2_X1 g_g7450 (g6090, g7195, g7450);
OR2_X1 g_g7575 (g7323, g7142, g7575);
OR2_X1 g_g7682 (g6044, g7412, g7682);
OR2_X1 g_g7687 (g6053, g7416, g7687);
OR2_X1 g_g7690 (g4181, g7417, g7690);
OR2_X1 g_g7697 (g7419, g3187, g7697);
OR2_X1 g_g7782 (g4783, g7598, g7782);
OR2_X1 g_g7783 (g4787, g7600, g7783);
OR3_X1 g_I14219 (g979, g7566, g1865, I14219);
OR4_X1 g_g7784 (g7406, g6664, g3492, I14219, g7784);
OR2_X1 g_g7787 (g4791, g7602, g7787);
OR2_X1 g_g7788 (g4794, g7604, g7788);
OR2_X1 g_g7791 (g4796, g7606, g7791);
OR2_X1 g_g7810 (g4799, g7609, g7810);
OR2_X1 g_g7825 (g4801, g7615, g7825);
OR2_X1 g_g7826 (g4804, g7626, g7826);
OR2_X1 g_g7834 (g7724, g6762, g7834);
OR3_X1 g_I14302 (g6664, g3492, g979, I14302);
OR4_X1 g_g8009 (g3591, g7406, g7566, I14302, g8009);
OR3_X1 g_g8082 (g7654, g7628, g7611, g8082);
OR3_X1 g_I14366 (g7566, g1030, g6664, I14366);
OR3_X1 g_g8091 (g7215, g6452, I14366, g8091);
OR3_X1 g_g8128 (g7566, g6910, g6452, g8128);
OR2_X1 g_g8146 (g6045, g7597, g8146);
OR2_X1 g_g8154 (g6054, g7607, g8154);
OR2_X1 g_g8155 (g7632, g3219, g8155);
OR4_X1 g_g8176 (g7566, g1030, g6664, g6452, g8176);
OR4_X1 g_I14467 (g7993, g7966, g7793, g7811, I14467);
OR4_X1 g_I14468 (g7937, g7887, g8029, g8018, I14468);
OR4_X1 g_I14479 (g7993, g7966, g7793, g7811, I14479);
OR4_X1 g_I14480 (g7937, g7887, g8029, g8018, I14480);
OR4_X1 g_I14484 (g7993, g7966, g7793, g7811, I14484);
OR4_X1 g_I14485 (g7937, g7887, g8029, g8018, I14485);
OR4_X1 g_I14495 (g7993, g7966, g7793, g7811, I14495);
OR4_X1 g_I14496 (g7937, g7887, g8029, g8018, I14496);
OR2_X1 g_g8613 (g8082, g7616, g8613);
OR2_X1 g_g8634 (g6047, g8060, g8634);
OR2_X1 g_g8637 (g6057, g8071, g8637);
OR4_X1 g_I14753 (g7993, g7966, g7793, g7811, I14753);
OR4_X1 g_I14754 (g7937, g7887, g8029, g8018, I14754);
OR4_X1 g_I14758 (g7993, g7966, g7793, g7811, I14758);
OR4_X1 g_I14759 (g7937, g7887, g8029, g8018, I14759);
OR4_X1 g_I14766 (g7993, g7966, g7793, g7811, I14766);
OR4_X1 g_I14767 (g7937, g7887, g8029, g8018, I14767);
OR4_X1 g_I14771 (g7993, g7966, g7793, g7811, I14771);
OR4_X1 g_I14772 (g7937, g7887, g8029, g8018, I14772);
OR3_X1 g_I14831 (g8483, g8464, g8514, I14831);
OR3_X1 g_I14834 (g8483, g8464, g8514, I14834);
OR4_X1 g_I14932 (g8278, g8329, g8461, g8382, I14932);
OR4_X1 g_I14933 (g8385, g8404, g8441, g8462, I14933);
OR3_X1 g_g8758 (g8655, I14932, I14933, g8758);
OR4_X1 g_I14941 (g8275, g8323, g8459, g8380, I14941);
OR4_X1 g_I14942 (g8439, g8440, g8405, g8460, I14942);
OR3_X1 g_g8763 (g8232, I14941, I14942, g8763);
OR4_X1 g_I14951 (g8328, g8316, g8455, g8378, I14951);
OR4_X1 g_I14952 (g8456, g8513, g8458, g8236, I14952);
OR2_X1 g_g8769 (I14951, I14952, g8769);
OR4_X1 g_I14959 (g8322, g8308, g8438, g8612, I14959);
OR4_X1 g_I14960 (g8621, g8622, g8628, g8230, I14960);
OR2_X1 g_g8773 (I14959, I14960, g8773);
OR4_X1 g_I14969 (g8315, g8377, g8359, g8611, I14969);
OR4_X1 g_I14970 (g8457, g8383, g8626, g8233, I14970);
OR2_X1 g_g8777 (I14969, I14970, g8777);
OR3_X1 g_I14980 (g8362, g8403, g8610, I14980);
OR3_X1 g_g8782 (g8624, g8659, I14980, g8782);
OR3_X1 g_I14985 (g8341, g8384, g8542, I14985);
OR3_X1 g_g8785 (g8623, g8656, I14985, g8785);
OR3_X1 g_I14990 (g8337, g8379, g8543, I14990);
OR3_X1 g_g8788 (g8620, g8658, I14990, g8788);
OR4_X1 g_g8794 (g8153, g8074, g8069, g8523, g8794);
OR4_X1 g_g8795 (g8151, g8077, g8075, g8279, g8795);
OR4_X1 g_g8796 (g8150, g8078, g8070, g8360, g8796);
OR4_X1 g_I15017 (g8131, g8111, g8042, g8156, I15017);
OR4_X1 g_I15018 (g7855, g7838, g7905, g7870, I15018);
OR4_X1 g_I15019 (g7951, g7920, g7983, g8181, I15019);
OR4_X1 g_I15020 (g8363, g8342, g8407, g8386, I15020);
OR4_X1 g_I15021 (I15017, I15018, I15019, I15020, I15021);
OR2_X1 g_g8804 (g6060, g8609, g8804);
OR4_X1 g_I15029 (g8131, g8111, g8042, g8156, I15029);
OR4_X1 g_I15030 (g7855, g7838, g7905, g7870, I15030);
OR4_X1 g_I15031 (g7951, g7920, g7983, g8181, I15031);
OR4_X1 g_I15032 (g8363, g8342, g8407, g8386, I15032);
OR4_X1 g_I15033 (I15029, I15030, I15031, I15032, I15033);
OR4_X1 g_I15040 (g8131, g8111, g8042, g8156, I15040);
OR4_X1 g_I15041 (g7855, g7838, g7905, g7870, I15041);
OR4_X1 g_I15042 (g7951, g7920, g7983, g8181, I15042);
OR4_X1 g_I15043 (g8363, g8342, g8407, g8386, I15043);
OR4_X1 g_I15044 (I15040, I15041, I15042, I15043, I15044);
OR4_X1 g_I15051 (g8131, g8111, g8042, g8156, I15051);
OR4_X1 g_I15052 (g7855, g7838, g7905, g7870, I15052);
OR4_X1 g_I15053 (g7951, g7920, g7983, g8181, I15053);
OR4_X1 g_I15054 (g8363, g8342, g8407, g8386, I15054);
OR4_X1 g_I15055 (I15051, I15052, I15053, I15054, I15055);
OR4_X1 g_I15071 (g8131, g8111, g8042, g8156, I15071);
OR4_X1 g_I15072 (g7855, g7838, g7905, g7870, I15072);
OR4_X1 g_I15073 (g7951, g7920, g7983, g8181, I15073);
OR4_X1 g_I15074 (g8363, g8342, g8407, g8386, I15074);
OR4_X1 g_I15075 (I15071, I15072, I15073, I15074, I15075);
OR4_X1 g_I15082 (g8131, g8111, g8042, g8156, I15082);
OR4_X1 g_I15083 (g7855, g7838, g7905, g7870, I15083);
OR4_X1 g_I15084 (g7951, g7920, g7983, g8181, I15084);
OR4_X1 g_I15085 (g8363, g8342, g8407, g8386, I15085);
OR4_X1 g_I15086 (I15082, I15083, I15084, I15085, I15086);
OR4_X1 g_I15098 (g8131, g8111, g8042, g8156, I15098);
OR4_X1 g_I15099 (g7855, g7838, g7905, g7870, I15099);
OR4_X1 g_I15100 (g7951, g7920, g7983, g8181, I15100);
OR4_X1 g_I15101 (g8363, g8342, g8407, g8386, I15101);
OR4_X1 g_I15102 (I15098, I15099, I15100, I15101, I15102);
OR4_X1 g_I15109 (g8131, g8111, g8042, g8156, I15109);
OR4_X1 g_I15110 (g7855, g7838, g7905, g7870, I15110);
OR4_X1 g_I15111 (g7951, g7920, g7983, g8181, I15111);
OR4_X1 g_I15112 (g8363, g8342, g8407, g8386, I15112);
OR4_X1 g_I15113 (I15109, I15110, I15111, I15112, I15113);
OR2_X1 g_g8834 (g7096, g8229, g8834);
OR3_X1 g_I15147 (g8483, g8464, g8514, I15147);
OR3_X1 g_I15152 (g8483, g8464, g8514, I15152);
OR3_X1 g_I15165 (g8483, g8464, g8514, I15165);
OR3_X1 g_I15169 (g8483, g8464, g8514, I15169);
OR3_X1 g_I15172 (g8483, g8464, g8514, I15172);
OR3_X1 g_I15175 (g8483, g8464, g8514, I15175);
OR4_X1 g_I15228 (g8270, g8258, g8281, g8273, I15228);
OR4_X1 g_I15229 (g8262, g8303, g8268, g8312, I15229);
OR4_X1 g_I15230 (g8274, g8321, g8298, g8696, I15230);
OR4_X1 g_I15231 (g8701, g8715, g8730, g8720, I15231);
OR4_X1 g_I15232 (I15228, I15229, I15230, I15231, I15232);
OR3_X1 g_g8884 (g8735, g8818, I15232, g8884);
OR4_X1 g_I15239 (g8264, g8260, g8277, g8301, I15239);
OR4_X1 g_I15240 (g8259, g8294, g8263, g8305, I15240);
OR4_X1 g_I15241 (g8269, g8314, g8309, g8695, I15241);
OR4_X1 g_I15242 (g8697, g8714, g8718, g8719, I15242);
OR4_X1 g_I15243 (I15239, I15240, I15241, I15242, I15243);
OR3_X1 g_g8885 (g8723, g8806, I15243, g8885);
OR4_X1 g_I15250 (g8238, g8265, g8272, g8292, I15250);
OR4_X1 g_I15251 (g8302, g8288, g8311, g8296, I15251);
OR4_X1 g_I15252 (g8320, g8307, g8317, g8692, I15252);
OR4_X1 g_I15253 (g8698, g8711, g8722, g8716, I15253);
OR4_X1 g_I15254 (I15250, I15251, I15252, I15253, I15254);
OR3_X1 g_g8886 (g8727, g8812, I15254, g8886);
OR4_X1 g_I15261 (g8256, g8271, g8267, g8286, I15261);
OR4_X1 g_I15262 (g8293, g8283, g8304, g8289, I15262);
OR4_X1 g_I15263 (g8313, g8297, g8310, g8690, I15263);
OR4_X1 g_I15264 (g8700, g8708, g8726, g8731, I15264);
OR4_X1 g_I15265 (I15261, I15262, I15263, I15264, I15265);
OR2_X1 g_g8887 (I15265, g8819, g8887);
OR4_X1 g_I15272 (g8237, g8300, g8261, g8282, I15272);
OR4_X1 g_I15273 (g8287, g8334, g8295, g8339, I15273);
OR4_X1 g_I15274 (g8306, g8361, g8299, g8687, I15274);
OR4_X1 g_I15275 (g8693, g8703, g8712, g8717, I15275);
OR4_X1 g_I15276 (I15272, I15273, I15274, I15275, I15276);
OR2_X1 g_g8888 (I15276, g8807, g8888);
OR4_X1 g_I15283 (g8291, g8276, g8325, g8330, I15283);
OR4_X1 g_I15284 (g8335, g8340, g8290, g8691, I15284);
OR3_X1 g_I15285 (g8709, g8713, g8803, I15285);
OR3_X1 g_g8889 (I15283, I15284, I15285, g8889);
OR4_X1 g_I15290 (g8285, g8266, g8318, g8326, I15290);
OR4_X1 g_I15291 (g8331, g8336, g8338, g8688, I15291);
OR3_X1 g_I15292 (g8704, g8710, g8805, I15292);
OR3_X1 g_g8890 (I15290, I15291, I15292, g8890);
OR4_X1 g_I15297 (g8280, g8257, g8319, g8327, I15297);
OR4_X1 g_I15298 (g8332, g8333, g8686, g8702, I15298);
OR4_X1 g_g8891 (g8705, g8811, I15297, I15298, g8891);
OR2_X1 g_g8893 (g8814, g8643, g8893);
OR2_X1 g_g8894 (g8817, g8645, g8894);
OR2_X1 g_g8895 (g8823, g8646, g8895);
OR2_X1 g_g8896 (g8828, g8648, g8896);
OR2_X1 g_g8897 (g8833, g8650, g8897);
OR2_X1 g_g8899 (g8839, g8652, g8899);
OR2_X1 g_g8900 (g8840, g8653, g8900);
OR2_X1 g_g8902 (g8844, g8654, g8902);
OR3_X1 g_g8904 (g8090, g8080, g8706, g8904);
OR3_X1 g_g8905 (g8089, g8087, g8694, g8905);
OR3_X1 g_g8906 (g8088, g8062, g8699, g8906);
OR3_X1 g_g8907 (g8081, g8064, g8707, g8907);
OR3_X1 g_g8908 (g8079, g8066, g8855, g8908);
OR2_X1 g_g8909 (g6043, g8764, g8909);
OR3_X1 g_I15400 (g8736, g8748, g8740, I15400);
OR3_X1 g_g8964 (g8915, g8863, I15400, g8964);
OR4_X1 g_g8965 (g8739, g8742, g8914, g8847, g8965);
OR4_X1 g_g8966 (g8741, g8745, g8912, g8850, g8966);
OR2_X1 g_g8979 (g8919, g8813, g8979);
OR2_X1 g_g8980 (g8920, g8815, g8980);
OR2_X1 g_g8981 (g8921, g8816, g8981);
OR2_X1 g_g8982 (g8922, g8820, g8982);
OR2_X1 g_g8983 (g8923, g8821, g8983);
OR2_X1 g_g8984 (g8924, g8822, g8984);
OR2_X1 g_g8985 (g8925, g8824, g8985);
OR2_X1 g_g8986 (g8926, g8825, g8986);
OR2_X1 g_g8987 (g8927, g8826, g8987);
OR2_X1 g_g8988 (g8928, g8827, g8988);
OR2_X1 g_g8989 (g8929, g8829, g8989);
OR2_X1 g_g8990 (g8930, g8830, g8990);
OR2_X1 g_g8991 (g8931, g8831, g8991);
OR2_X1 g_g8992 (g8932, g8832, g8992);
OR2_X1 g_g8993 (g8933, g8835, g8993);
OR2_X1 g_g8994 (g8934, g8836, g8994);
OR2_X1 g_g8995 (g8935, g8837, g8995);
OR2_X1 g_g8996 (g8936, g8838, g8996);
OR2_X1 g_g8997 (g8937, g8841, g8997);
OR2_X1 g_g8998 (g8938, g8842, g8998);
OR2_X1 g_g8999 (g8939, g8843, g8999);
OR2_X1 g_g9000 (g8940, g8845, g9000);
OR2_X1 g_g9001 (g8941, g8846, g9001);
OR2_X1 g_g9002 (g8942, g8848, g9002);
OR2_X1 g_g9003 (g8943, g8849, g9003);
OR2_X1 g_g9004 (g8944, g8851, g9004);
OR2_X1 g_g9005 (g8945, g8852, g9005);
OR2_X1 g_g9006 (g8946, g8853, g9006);
OR2_X1 g_g9007 (g8947, g8854, g9007);
OR2_X1 g_g9008 (g8948, g8857, g9008);
OR2_X1 g_g9009 (g8949, g8858, g9009);
OR2_X1 g_g9010 (g8950, g8860, g9010);
OR2_X1 g_g9011 (g6046, g8892, g9011);
OR4_X1 g_g9046 (g8744, g8749, g9016, g8862, g9046);
OR4_X1 g_g9049 (g8732, g8737, g9015, g8861, g9049);
OR4_X1 g_g9052 (g8728, g8733, g9014, g8679, g9052);
OR4_X1 g_g9054 (g8724, g8729, g9013, g8680, g9054);
OR4_X1 g_g9055 (g8721, g8725, g9012, g8859, g9055);
OR2_X1 g_g9122 (g8953, g9084, g9122);
OR2_X1 g_g9123 (g8954, g9037, g9123);
OR2_X1 g_g9124 (g8876, g9038, g9124);
OR2_X1 g_g9135 (g8951, g9130, g9135);
OR2_X1 g_g9136 (g8952, g9131, g9136);
OR2_X1 g_g9137 (g8877, g9118, g9137);
OR2_X1 g_g9138 (g8878, g9119, g9138);
OR2_X1 g_g9139 (g8879, g9120, g9139);
OR2_X1 g_g9148 (g9143, g9024, g9148);
OR2_X1 g_g9151 (g9144, g8961, g9151);
OR2_X1 g_g9154 (g9142, g9021, g9154);
OR2_X1 g_g9162 (g9158, g9022, g9162);
OR2_X1 g_g9165 (g9159, g9023, g9165);
OR2_X1 g_g9168 (g9160, g9025, g9168);
OR2_X1 g_g9171 (g9146, g8962, g9171);
OR2_X1 g_g9174 (g9147, g8963, g9174);
OR2_X1 g_g9239 (g7653, g9226, g9239);
OR2_X1 g_g9261 (g9238, g6227, g9261);
OR2_X1 g_g9264 (g9247, g6242, g9264);
OR2_X1 g_g9267 (g9251, g6225, g9267);
OR2_X1 g_g9282 (g9270, g6238, g9282);
OR2_X1 g_g9285 (g9271, g6221, g9285);
OR2_X1 g_g9288 (g9272, g6235, g9288);
OR2_X1 g_g9291 (g9273, g6216, g9291);
OR2_X1 g_g9294 (g9274, g6230, g9294);
OR2_X1 g_g9337 (g9240, g9327, g9337);
OR2_X1 g_g9338 (g9258, g9334, g9338);
OR2_X1 g_g9339 (g9259, g9335, g9339);
OR2_X1 g_g9352 (g9343, g4526, g9352);
OR2_X1 g_g9354 (g9275, g9344, g9354);
OR2_X1 g_g9355 (g9276, g9345, g9355);
OR2_X1 g_g9356 (g9277, g9346, g9356);
OR2_X1 g_g9357 (g9278, g9347, g9357);
OR2_X1 g_g9358 (g9279, g9348, g9358);
OR2_X1 g_g9363 (g9359, g6210, g9363);
OR2_X1 g_g9377 (g9371, g6757, g9377);
OR2_X1 g_g9387 (g9349, g9384, g9387);
NAND2_X1 g_I5505 (g1532, g1528, I5505);
NAND2_X1 g_I5506 (g1532, I5505, I5506);
NAND2_X1 g_I5507 (g1528, I5505, I5507);
NAND2_X1 g_g1678 (I5506, I5507, g1678);
NAND2_X1 g_I5519 (g1087, g1098, I5519);
NAND2_X1 g_I5520 (g1087, I5519, I5520);
NAND2_X1 g_I5521 (g1098, I5519, I5521);
NAND2_X1 g_g1682 (I5520, I5521, g1682);
NAND2_X1 g_I5598 (g1481, g1489, I5598);
NAND2_X1 g_I5599 (g1481, I5598, I5599);
NAND2_X1 g_I5600 (g1489, I5598, I5600);
NAND2_X1 g_g1759 (I5599, I5600, g1759);
NAND2_X1 g_I5619 (g1092, g1130, I5619);
NAND2_X1 g_I5620 (g1092, I5619, I5620);
NAND2_X1 g_I5621 (g1130, I5619, I5621);
NAND2_X1 g_g1775 (I5620, I5621, g1775);
NAND2_X1 g_I5695 (g1513, g1524, I5695);
NAND2_X1 g_I5696 (g1513, I5695, I5696);
NAND2_X1 g_I5697 (g1524, I5695, I5697);
NAND2_X1 g_g1819 (I5696, I5697, g1819);
NAND2_X1 g_g1910 (g1435, g1439, g1910);
NAND2_X1 g_g2051 (g1444, g1450, g2051);
NAND2_X1 g_I6064 (g852, g883, I6064);
NAND2_X1 g_I6065 (g852, I6064, I6065);
NAND2_X1 g_I6066 (g883, I6064, I6066);
NAND2_X1 g_g2294 (I6065, I6066, g2294);
NAND2_X1 g_I6102 (g849, g921, I6102);
NAND2_X1 g_I6103 (g849, I6102, I6103);
NAND2_X1 g_I6104 (g921, I6102, I6104);
NAND2_X1 g_g2315 (I6103, I6104, g2315);
NAND2_X1 g_I6133 (g846, g916, I6133);
NAND2_X1 g_I6134 (g846, I6133, I6134);
NAND2_X1 g_I6135 (g916, I6133, I6135);
NAND2_X1 g_g2330 (I6134, I6135, g2330);
NAND2_X1 g_g2333 (g985, g990, g2333);
NAND2_X1 g_I6170 (g843, g911, I6170);
NAND2_X1 g_I6171 (g843, I6170, I6171);
NAND2_X1 g_I6172 (g911, I6170, I6172);
NAND2_X1 g_g2352 (I6171, I6172, g2352);
NAND2_X1 g_I6201 (g831, g891, I6201);
NAND2_X1 g_I6202 (g831, I6201, I6202);
NAND2_X1 g_I6203 (g891, I6201, I6203);
NAND2_X1 g_g2367 (I6202, I6203, g2367);
NAND2_X1 g_I6232 (g834, g896, I6232);
NAND2_X1 g_I6233 (g834, I6232, I6233);
NAND2_X1 g_I6234 (g896, I6232, I6234);
NAND2_X1 g_g2378 (I6233, I6234, g2378);
NAND2_X1 g_I6257 (g837, g901, I6257);
NAND2_X1 g_I6258 (g837, I6257, I6258);
NAND2_X1 g_I6259 (g901, I6257, I6259);
NAND2_X1 g_g2385 (I6258, I6259, g2385);
NAND2_X1 g_I6273 (g840, g906, I6273);
NAND2_X1 g_I6274 (g840, I6273, I6274);
NAND2_X1 g_I6275 (g906, I6273, I6275);
NAND2_X1 g_g2395 (I6274, I6275, g2395);
NAND2_X1 g_g2474 (g1405, g1412, g2474);
NAND2_X1 g_I6499 (g1913, g1537, I6499);
NAND2_X1 g_I6500 (g1913, I6499, I6500);
NAND2_X1 g_I6501 (g1537, I6499, I6501);
NAND2_X1 g_g2751 (I6500, I6501, g2751);
NAND2_X1 g_I6522 (g1919, g1102, I6522);
NAND2_X1 g_I6523 (g1919, I6522, I6523);
NAND2_X1 g_I6524 (g1102, I6522, I6524);
NAND2_X1 g_g2783 (I6523, I6524, g2783);
NAND2_X1 g_I6538 (g2555, g2557, I6538);
NAND2_X1 g_I6539 (g2555, I6538, I6539);
NAND2_X1 g_I6540 (g2557, I6538, I6540);
NAND2_X1 g_g2801 (I6539, I6540, g2801);
NAND2_X1 g_I6739 (g195, g1970, I6739);
NAND2_X1 g_I6740 (g195, I6739, I6740);
NAND2_X1 g_I6741 (g1970, I6739, I6741);
NAND2_X1 g_g2995 (I6740, I6741, g2995);
NAND2_X1 g_I6750 (g1733, g1494, I6750);
NAND2_X1 g_I6751 (g1733, I6750, I6751);
NAND2_X1 g_I6752 (g1494, I6750, I6752);
NAND2_X1 g_g3011 (I6751, I6752, g3011);
NAND2_X1 g_I6757 (g186, g1983, I6757);
NAND2_X1 g_I6758 (g186, I6757, I6758);
NAND2_X1 g_I6759 (g1983, I6757, I6759);
NAND2_X1 g_g3012 (I6758, I6759, g3012);
NAND2_X1 g_I6774 (g2386, g1134, I6774);
NAND2_X1 g_I6775 (g2386, I6774, I6775);
NAND2_X1 g_I6776 (g1134, I6774, I6776);
NAND2_X1 g_g3028 (I6775, I6776, g3028);
NAND2_X1 g_I6813 (g210, g2052, I6813);
NAND2_X1 g_I6814 (g210, I6813, I6814);
NAND2_X1 g_I6815 (g2052, I6813, I6815);
NAND2_X1 g_g3083 (I6814, I6815, g3083);
NAND2_X1 g_I6842 (g205, g2016, I6842);
NAND2_X1 g_I6843 (g205, I6842, I6843);
NAND2_X1 g_I6844 (g2016, I6842, I6844);
NAND2_X1 g_g3129 (I6843, I6844, g3129);
NAND2_X1 g_I6876 (g1967, g1910, I6876);
NAND2_X1 g_I6877 (g1967, I6876, I6877);
NAND2_X1 g_I6878 (g1910, I6876, I6878);
NAND2_X1 g_g3221 (I6877, I6878, g3221);
NAND2_X1 g_g3231 (g1889, g1904, g3231);
NAND2_X1 g_g3232 (g2298, g2276, g3232);
NAND2_X1 g_I6904 (g2105, g1838, I6904);
NAND2_X1 g_I6905 (g2105, I6904, I6905);
NAND2_X1 g_I6906 (g1838, I6904, I6906);
NAND2_X1 g_g3286 (I6905, I6906, g3286);
NAND2_X1 g_I6916 (g2360, g1732, I6916);
NAND2_X1 g_I6917 (g2360, I6916, I6917);
NAND2_X1 g_I6918 (g1732, I6916, I6918);
NAND2_X1 g_g3314 (I6917, I6918, g3314);
NAND2_X1 g_I6923 (g1728, g33, I6923);
NAND2_X1 g_I6924 (g1728, I6923, I6924);
NAND2_X1 g_I6925 (g33, I6923, I6925);
NAND2_X1 g_g3315 (I6924, I6925, g3315);
NAND2_X1 g_I6939 (g2161, g2051, I6939);
NAND2_X1 g_I6940 (g2161, I6939, I6940);
NAND2_X1 g_I6941 (g2051, I6939, I6941);
NAND2_X1 g_g3358 (I6940, I6941, g3358);
NAND2_X1 g_I6996 (g2275, g2242, I6996);
NAND2_X1 g_I6997 (g2275, I6996, I6997);
NAND2_X1 g_I6998 (g2242, I6996, I6998);
NAND2_X1 g_g3518 (I6997, I6998, g3518);
NAND2_X1 g_I7009 (g2295, g2333, I7009);
NAND2_X1 g_I7010 (g2295, I7009, I7010);
NAND2_X1 g_I7011 (g2333, I7009, I7011);
NAND2_X1 g_g3525 (I7010, I7011, g3525);
NAND2_X1 g_I7068 (g1639, g1643, I7068);
NAND2_X1 g_I7069 (g1639, I7068, I7069);
NAND2_X1 g_I7070 (g1643, I7068, I7070);
NAND2_X1 g_g3602 (I7069, I7070, g3602);
NAND2_X1 g_I7085 (g1753, g1918, I7085);
NAND2_X1 g_I7086 (g1753, I7085, I7086);
NAND2_X1 g_I7087 (g1918, I7085, I7087);
NAND2_X1 g_g3613 (I7086, I7087, g3613);
NAND2_X1 g_I7138 (g2404, g2397, I7138);
NAND2_X1 g_I7139 (g2404, I7138, I7139);
NAND2_X1 g_I7140 (g2397, I7138, I7140);
NAND2_X1 g_g3656 (I7139, I7140, g3656);
NAND2_X1 g_I7148 (g799, g1974, I7148);
NAND2_X1 g_I7149 (g799, I7148, I7149);
NAND2_X1 g_I7150 (g1974, I7148, I7150);
NAND2_X1 g_g3658 (I7149, I7150, g3658);
NAND2_X1 g_I7156 (g2331, g929, I7156);
NAND2_X1 g_I7157 (g2331, I7156, I7157);
NAND2_X1 g_I7158 (g929, I7156, I7158);
NAND2_X1 g_g3665 (I7157, I7158, g3665);
NAND2_X1 g_I7172 (g1739, g2006, I7172);
NAND2_X1 g_I7173 (g1739, I7172, I7173);
NAND2_X1 g_I7174 (g2006, I7172, I7174);
NAND2_X1 g_g3678 (I7173, I7174, g3678);
NAND2_X1 g_I7179 (g2351, g795, I7179);
NAND2_X1 g_I7180 (g2351, I7179, I7180);
NAND2_X1 g_I7181 (g795, I7179, I7181);
NAND2_X1 g_g3679 (I7180, I7181, g3679);
NAND2_X1 g_I7186 (g2353, g1834, I7186);
NAND2_X1 g_I7187 (g2353, I7186, I7187);
NAND2_X1 g_I7188 (g1834, I7186, I7188);
NAND2_X1 g_g3680 (I7187, I7188, g3680);
NAND2_X1 g_g3681 (g866, g2368, g3681);
NAND2_X1 g_g3706 (g1556, g2510, g3706);
NAND2_X1 g_I7214 (g815, g2091, I7214);
NAND2_X1 g_I7215 (g815, I7214, I7215);
NAND2_X1 g_I7216 (g2091, I7214, I7216);
NAND2_X1 g_g3722 (I7215, I7216, g3722);
NAND2_X1 g_I7239 (g1658, g2134, I7239);
NAND2_X1 g_I7240 (g1658, I7239, I7240);
NAND2_X1 g_I7241 (g2134, I7239, I7241);
NAND2_X1 g_g3767 (I7240, I7241, g3767);
NAND2_X1 g_I7268 (g2486, g955, I7268);
NAND2_X1 g_I7269 (g2486, I7268, I7269);
NAND2_X1 g_I7270 (g955, I7268, I7270);
NAND2_X1 g_g3811 (I7269, I7270, g3811);
NAND2_X1 g_I7277 (g2497, g1898, I7277);
NAND2_X1 g_I7278 (g2497, I7277, I7278);
NAND2_X1 g_I7279 (g1898, I7277, I7279);
NAND2_X1 g_g3818 (I7278, I7279, g3818);
NAND2_X1 g_g3883 (g2276, g3188, g3883);
NAND2_X1 g_I7421 (g2525, g2703, I7421);
NAND2_X1 g_I7422 (g2525, I7421, I7422);
NAND2_X1 g_I7423 (g2703, I7421, I7423);
NAND2_X1 g_g3886 (I7422, I7423, g3886);
NAND2_X1 g_I7428 (g3222, g1541, I7428);
NAND2_X1 g_I7429 (g3222, I7428, I7429);
NAND2_X1 g_I7430 (g1541, I7428, I7430);
NAND2_X1 g_g3887 (I7429, I7430, g3887);
NAND2_X1 g_I7436 (g2517, g3822, I7436);
NAND2_X1 g_I7437 (g2517, I7436, I7437);
NAND2_X1 g_I7438 (g3822, I7436, I7438);
NAND2_X1 g_g3889 (I7437, I7438, g3889);
NAND2_X1 g_I7443 (g2973, g1701, I7443);
NAND2_X1 g_I7444 (g2973, I7443, I7444);
NAND2_X1 g_I7445 (g1701, I7443, I7445);
NAND2_X1 g_g3890 (I7444, I7445, g3890);
NAND2_X1 g_I7452 (g3226, g1106, I7452);
NAND2_X1 g_I7453 (g3226, I7452, I7453);
NAND2_X1 g_I7454 (g1106, I7452, I7454);
NAND2_X1 g_g3893 (I7453, I7454, g3893);
NAND2_X1 g_I7459 (g2506, g3815, I7459);
NAND2_X1 g_I7460 (g2506, I7459, I7460);
NAND2_X1 g_I7461 (g3815, I7459, I7461);
NAND2_X1 g_g3894 (I7460, I7461, g3894);
NAND2_X1 g_I7466 (g2982, g1704, I7466);
NAND2_X1 g_I7467 (g2982, I7466, I7467);
NAND2_X1 g_I7468 (g1704, I7466, I7468);
NAND2_X1 g_g3895 (I7467, I7468, g3895);
NAND2_X1 g_I7478 (g2502, g3808, I7478);
NAND2_X1 g_I7479 (g2502, I7478, I7479);
NAND2_X1 g_I7480 (g3808, I7478, I7480);
NAND2_X1 g_g3899 (I7479, I7480, g3899);
NAND2_X1 g_I7485 (g2989, g1708, I7485);
NAND2_X1 g_I7486 (g2989, I7485, I7486);
NAND2_X1 g_I7487 (g1708, I7485, I7487);
NAND2_X1 g_g3900 (I7486, I7487, g3900);
NAND2_X1 g_I7503 (g2498, g3802, I7503);
NAND2_X1 g_I7504 (g2498, I7503, I7504);
NAND2_X1 g_I7505 (g3802, I7503, I7505);
NAND2_X1 g_g3906 (I7504, I7505, g3906);
NAND2_X1 g_I7510 (g2992, g1711, I7510);
NAND2_X1 g_I7511 (g2992, I7510, I7511);
NAND2_X1 g_I7512 (g1711, I7510, I7512);
NAND2_X1 g_g3907 (I7511, I7512, g3907);
NAND2_X1 g_I7531 (g2487, g3787, I7531);
NAND2_X1 g_I7532 (g2487, I7531, I7532);
NAND2_X1 g_I7533 (g3787, I7531, I7533);
NAND2_X1 g_g3914 (I7532, I7533, g3914);
NAND2_X1 g_I7538 (g2996, g1715, I7538);
NAND2_X1 g_I7539 (g2996, I7538, I7539);
NAND2_X1 g_I7540 (g1715, I7538, I7540);
NAND2_X1 g_g3915 (I7539, I7540, g3915);
NAND2_X1 g_I7567 (g2481, g3780, I7567);
NAND2_X1 g_I7568 (g2481, I7567, I7568);
NAND2_X1 g_I7569 (g3780, I7567, I7569);
NAND2_X1 g_g3924 (I7568, I7569, g3924);
NAND2_X1 g_I7574 (g2999, g1718, I7574);
NAND2_X1 g_I7575 (g2999, I7574, I7575);
NAND2_X1 g_I7576 (g1718, I7574, I7576);
NAND2_X1 g_g3925 (I7575, I7576, g3925);
NAND2_X1 g_I7609 (g2471, g3771, I7609);
NAND2_X1 g_I7610 (g2471, I7609, I7610);
NAND2_X1 g_I7611 (g3771, I7609, I7611);
NAND2_X1 g_g3938 (I7610, I7611, g3938);
NAND2_X1 g_I7616 (g3008, g1721, I7616);
NAND2_X1 g_I7617 (g3008, I7616, I7617);
NAND2_X1 g_I7618 (g1721, I7616, I7618);
NAND2_X1 g_g3939 (I7617, I7618, g3939);
NAND2_X1 g_I7891 (g2979, g1499, I7891);
NAND2_X1 g_I7892 (g2979, I7891, I7892);
NAND2_X1 g_I7893 (g1499, I7891, I7893);
NAND2_X1 g_g4090 (I7892, I7893, g4090);
NAND2_X1 g_I7937 (g3614, g1138, I7937);
NAND2_X1 g_I7938 (g3614, I7937, I7938);
NAND2_X1 g_I7939 (g1138, I7937, I7939);
NAND2_X1 g_g4110 (I7938, I7939, g4110);
NAND2_X1 g_I8119 (g1904, g3220, I8119);
NAND2_X1 g_I8120 (g1904, I8119, I8120);
NAND2_X1 g_I8121 (g3220, I8119, I8121);
NAND2_X1 g_g4219 (I8120, I8121, g4219);
NAND2_X1 g_I8132 (g3232, g1646, I8132);
NAND2_X1 g_I8133 (g3232, I8132, I8133);
NAND2_X1 g_I8134 (g1646, I8132, I8134);
NAND2_X1 g_g4227 (I8133, I8134, g4227);
NAND2_X1 g_g4228 (g1408, g2665, g4228);
NAND2_X1 g_g4231 (g2276, g3258, g4231);
NAND2_X1 g_g4235 (g1415, g2668, g4235);
NAND2_X1 g_I8150 (g3229, g38, I8150);
NAND2_X1 g_I8151 (g3229, I8150, I8151);
NAND2_X1 g_I8152 (g38, I8150, I8152);
NAND2_X1 g_g4237 (I8151, I8152, g4237);
NAND2_X1 g_I8164 (g1943, g3231, I8164);
NAND2_X1 g_I8165 (g1943, I8164, I8165);
NAND2_X1 g_I8166 (g3231, I8164, I8166);
NAND2_X1 g_g4243 (I8165, I8166, g4243);
NAND2_X1 g_g4244 (g3549, g3533, g4244);
NAND2_X1 g_g4252 (g2276, g3313, g4252);
NAND2_X1 g_g4256 (g3233, g1444, g4256);
NAND2_X1 g_g4263 (g3260, g1435, g4263);
NAND2_X1 g_I8243 (g2011, g3506, I8243);
NAND2_X1 g_I8244 (g2011, I8243, I8244);
NAND2_X1 g_I8245 (g3506, I8243, I8245);
NAND2_X1 g_g4294 (I8244, I8245, g4294);
NAND2_X1 g_I8253 (g2454, g3825, I8253);
NAND2_X1 g_I8254 (g2454, I8253, I8254);
NAND2_X1 g_I8255 (g3825, I8253, I8255);
NAND2_X1 g_g4298 (I8254, I8255, g4298);
NAND3_X1 g_g4305 (g3712, g3700, g3732, g4305);
NAND3_X1 g_g4309 (g3002, g3124, g3659, g4309);
NAND2_X1 g_g4310 (g3666, g2460, g4310);
NAND2_X1 g_g4313 (g3712, g3700, g4313);
NAND2_X1 g_g4332 (g3681, g2368, g4332);
NAND2_X1 g_I8326 (g2011, g2721, I8326);
NAND2_X1 g_I8327 (g2011, I8326, I8327);
NAND2_X1 g_I8328 (g2721, I8326, I8328);
NAND2_X1 g_g4359 (I8327, I8328, g4359);
NAND2_X1 g_I8338 (g2966, g1698, I8338);
NAND2_X1 g_I8339 (g2966, I8338, I8339);
NAND2_X1 g_I8340 (g1698, I8338, I8340);
NAND2_X1 g_g4363 (I8339, I8340, g4363);
NAND2_X1 g_I8392 (g2949, g1925, I8392);
NAND2_X1 g_I8393 (g2949, I8392, I8393);
NAND2_X1 g_I8394 (g1925, I8392, I8394);
NAND2_X1 g_g4399 (I8393, I8394, g4399);
NAND2_X1 g_I8470 (g2525, g2821, I8470);
NAND2_X1 g_I8471 (g2525, I8470, I8471);
NAND2_X1 g_I8472 (g2821, I8470, I8472);
NAND2_X1 g_g4456 (I8471, I8472, g4456);
NAND2_X1 g_I8502 (g2986, g2038, I8502);
NAND2_X1 g_I8503 (g2986, I8502, I8503);
NAND2_X1 g_I8504 (g2038, I8502, I8504);
NAND2_X1 g_g4474 (I8503, I8504, g4474);
NAND2_X1 g_I8510 (g2517, g2807, I8510);
NAND2_X1 g_I8511 (g2517, I8510, I8511);
NAND2_X1 g_I8512 (g2807, I8510, I8512);
NAND2_X1 g_g4476 (I8511, I8512, g4476);
NAND2_X1 g_I8536 (g2506, g2798, I8536);
NAND2_X1 g_I8537 (g2506, I8536, I8537);
NAND2_X1 g_I8538 (g2798, I8536, I8538);
NAND2_X1 g_g4492 (I8537, I8538, g4492);
NAND2_X1 g_I8558 (g2502, g2790, I8558);
NAND2_X1 g_I8559 (g2502, I8558, I8559);
NAND2_X1 g_I8560 (g2790, I8558, I8560);
NAND2_X1 g_g4502 (I8559, I8560, g4502);
NAND2_X1 g_I8581 (g2498, g2777, I8581);
NAND2_X1 g_I8582 (g2498, I8581, I8582);
NAND2_X1 g_I8583 (g2777, I8581, I8583);
NAND2_X1 g_g4513 (I8582, I8583, g4513);
NAND2_X1 g_I8605 (g2487, g2764, I8605);
NAND2_X1 g_I8606 (g2487, I8605, I8606);
NAND2_X1 g_I8607 (g2764, I8605, I8607);
NAND2_X1 g_g4528 (I8606, I8607, g4528);
NAND2_X1 g_I8635 (g2481, g2743, I8635);
NAND2_X1 g_I8636 (g2481, I8635, I8636);
NAND2_X1 g_I8637 (g2743, I8635, I8637);
NAND2_X1 g_g4548 (I8636, I8637, g4548);
NAND2_X1 g_I8658 (g2471, g2724, I8658);
NAND2_X1 g_I8659 (g2471, I8658, I8659);
NAND2_X1 g_I8660 (g2724, I8658, I8660);
NAND2_X1 g_g4563 (I8659, I8660, g4563);
NAND2_X1 g_I8678 (g2467, g2706, I8678);
NAND2_X1 g_I8679 (g2467, I8678, I8679);
NAND2_X1 g_I8680 (g2706, I8678, I8680);
NAND2_X1 g_g4575 (I8679, I8680, g4575);
NAND2_X1 g_I8938 (g4239, g1545, I8938);
NAND2_X1 g_I8939 (g4239, I8938, I8939);
NAND2_X1 g_I8940 (g1545, I8938, I8940);
NAND2_X1 g_g4679 (I8939, I8940, g4679);
NAND2_X1 g_I8955 (g4246, g1110, I8955);
NAND2_X1 g_I8956 (g4246, I8955, I8956);
NAND2_X1 g_I8957 (g1110, I8955, I8957);
NAND2_X1 g_g4686 (I8956, I8957, g4686);
NAND2_X1 g_g4700 (g2460, g4271, g4700);
NAND3_X1 g_g4714 (g4344, g4335, g4328, g4714);
NAND2_X1 g_I9057 (g4059, g1504, I9057);
NAND2_X1 g_I9058 (g4059, I9057, I9058);
NAND2_X1 g_I9059 (g1504, I9057, I9059);
NAND2_X1 g_g4741 (I9058, I9059, g4741);
NAND2_X1 g_I9069 (g4400, g1149, I9069);
NAND2_X1 g_I9070 (g4400, I9069, I9070);
NAND2_X1 g_I9071 (g1149, I9069, I9071);
NAND2_X1 g_g4745 (I9070, I9071, g4745);
NAND2_X1 g_I9151 (g3883, g1649, I9151);
NAND2_X1 g_I9152 (g3883, I9151, I9152);
NAND2_X1 g_I9153 (g1649, I9151, I9153);
NAND2_X1 g_g4810 (I9152, I9153, g4810);
NAND2_X1 g_I9169 (g1935, g4244, I9169);
NAND2_X1 g_I9170 (g1935, I9169, I9170);
NAND2_X1 g_I9171 (g4244, I9169, I9171);
NAND2_X1 g_g4820 (I9170, I9171, g4820);
NAND2_X1 g_g4821 (g4220, g3605, g4821);
NAND2_X1 g_I9181 (g4231, g2007, I9181);
NAND2_X1 g_I9182 (g4231, I9181, I9182);
NAND2_X1 g_I9183 (g2007, I9181, I9183);
NAND2_X1 g_g4824 (I9182, I9183, g4824);
NAND3_X1 g_g4831 (g3635, g3605, g4220, g4831);
NAND2_X1 g_I9194 (g4252, g1652, I9194);
NAND2_X1 g_I9195 (g4252, I9194, I9195);
NAND2_X1 g_I9196 (g1652, I9194, I9196);
NAND2_X1 g_g4835 (I9195, I9196, g4835);
NAND2_X1 g_g4836 (g4288, g1879, g4836);
NAND2_X1 g_g4839 (g1879, g4269, g4839);
NAND2_X1 g_g4869 (g4254, g3533, g4869);
NAND4_X1 g_g4871 (g3635, g3605, g4220, g3644, g4871);
NAND4_X1 g_g4879 (g2595, g2584, g4270, g4281, g4879);
NAND2_X1 g_g4880 (g4287, g1879, g4880);
NAND2_X1 g_g4881 (g2460, g4315, g4881);
NAND2_X1 g_I9233 (g4310, g2180, I9233);
NAND2_X1 g_I9234 (g4310, I9233, I9234);
NAND2_X1 g_I9235 (g2180, I9233, I9235);
NAND2_X1 g_g4887 (I9234, I9235, g4887);
NAND2_X1 g_I9241 (g2540, g4305, I9241);
NAND2_X1 g_I9242 (g2540, I9241, I9242);
NAND2_X1 g_I9243 (g4305, I9241, I9243);
NAND2_X1 g_g4889 (I9242, I9243, g4889);
NAND2_X1 g_g4893 (g2460, g4312, g4893);
NAND2_X1 g_g4905 (g4282, g3533, g4905);
NAND2_X1 g_g4910 (g2460, g4314, g4910);
NAND2_X1 g_g4911 (g4320, g2044, g4911);
NAND2_X1 g_I9276 (g2533, g4313, I9276);
NAND2_X1 g_I9277 (g2533, I9276, I9277);
NAND2_X1 g_I9278 (g4313, I9276, I9278);
NAND2_X1 g_g4912 (I9277, I9278, g4912);
NAND2_X1 g_g4954 (g4319, g2460, g4954);
NAND2_X1 g_I9381 (g4062, g1908, I9381);
NAND2_X1 g_I9382 (g4062, I9381, I9382);
NAND2_X1 g_I9383 (g1908, I9381, I9383);
NAND2_X1 g_g5035 (I9382, I9383, g5035);
NAND2_X1 g_I9475 (g4038, g1942, I9475);
NAND2_X1 g_I9476 (g4038, I9475, I9476);
NAND2_X1 g_I9477 (g1942, I9475, I9477);
NAND2_X1 g_g5095 (I9476, I9477, g5095);
NAND2_X1 g_I9547 (g1952, g4307, I9547);
NAND2_X1 g_I9548 (g1952, I9547, I9548);
NAND2_X1 g_I9549 (g4307, I9547, I9549);
NAND2_X1 g_g5141 (I9548, I9549, g5141);
NAND2_X1 g_I9691 (g5096, g1037, I9691);
NAND2_X1 g_I9692 (g5096, I9691, I9692);
NAND2_X1 g_I9693 (g1037, I9691, I9693);
NAND2_X1 g_g5189 (I9692, I9693, g5189);
NAND2_X1 g_I9745 (g4826, g1549, I9745);
NAND2_X1 g_I9746 (g4826, I9745, I9746);
NAND2_X1 g_I9747 (g1549, I9745, I9747);
NAND2_X1 g_g5239 (I9746, I9747, g5239);
NAND2_X1 g_I9767 (g4832, g1114, I9767);
NAND2_X1 g_I9768 (g4832, I9767, I9768);
NAND2_X1 g_I9769 (g1114, I9767, I9769);
NAND2_X1 g_g5257 (I9768, I9769, g5257);
NAND3_X1 g_g5284 (g4344, g4335, g4963, g5284);
NAND3_X1 g_g5291 (g4344, g5002, g4963, g5291);
NAND3_X1 g_g5305 (g5009, g4335, g4328, g5305);
NAND3_X1 g_g5310 (g5009, g4335, g4963, g5310);
NAND3_X1 g_g5312 (g5009, g5002, g4963, g5312);
NAND2_X1 g_I9826 (g4729, g1509, I9826);
NAND2_X1 g_I9827 (g4729, I9826, I9827);
NAND2_X1 g_I9828 (g1509, I9826, I9828);
NAND2_X1 g_g5363 (I9827, I9828, g5363);
NAND2_X1 g_g5512 (g1879, g4877, g5512);
NAND2_X1 g_g5538 (g5132, g1266, g5538);
NAND2_X1 g_I9946 (g2128, g4905, I9946);
NAND2_X1 g_I9947 (g2128, I9946, I9947);
NAND2_X1 g_I9948 (g4905, I9946, I9948);
NAND2_X1 g_g5539 (I9947, I9948, g5539);
NAND2_X1 g_I9953 (g2131, g4831, I9953);
NAND2_X1 g_I9954 (g2131, I9953, I9954);
NAND2_X1 g_I9955 (g4831, I9953, I9955);
NAND2_X1 g_g5540 (I9954, I9955, g5540);
NAND2_X1 g_I9963 (g1938, g4869, I9963);
NAND2_X1 g_I9964 (g1938, I9963, I9964);
NAND2_X1 g_I9965 (g4869, I9963, I9965);
NAND2_X1 g_g5546 (I9964, I9965, g5546);
NAND2_X1 g_g5550 (g1879, g4830, g5550);
NAND2_X1 g_I9978 (g4880, g2092, I9978);
NAND2_X1 g_I9979 (g4880, I9978, I9979);
NAND2_X1 g_I9980 (g2092, I9978, I9980);
NAND2_X1 g_g5555 (I9979, I9980, g5555);
NAND2_X1 g_I9985 (g4836, g2096, I9985);
NAND2_X1 g_I9986 (g4836, I9985, I9986);
NAND2_X1 g_I9987 (g2096, I9985, I9987);
NAND2_X1 g_g5556 (I9986, I9987, g5556);
NAND2_X1 g_I9992 (g2145, g4871, I9992);
NAND2_X1 g_I9993 (g2145, I9992, I9993);
NAND2_X1 g_I9994 (g4871, I9992, I9994);
NAND2_X1 g_g5557 (I9993, I9994, g5557);
NAND2_X1 g_I9999 (g4839, g1929, I9999);
NAND2_X1 g_I10000 (g4839, I9999, I10000);
NAND2_X1 g_I10001 (g1929, I9999, I10001);
NAND2_X1 g_g5558 (I10000, I10001, g5558);
NAND2_X1 g_g5559 (g5132, g1257, g5559);
NAND2_X1 g_I10009 (g1949, g4821, I10009);
NAND2_X1 g_I10010 (g1949, I10009, I10010);
NAND2_X1 g_I10011 (g4821, I10009, I10011);
NAND2_X1 g_g5562 (I10010, I10011, g5562);
NAND2_X1 g_I10017 (g4700, g2174, I10017);
NAND2_X1 g_I10018 (g4700, I10017, I10018);
NAND2_X1 g_I10019 (g2174, I10017, I10019);
NAND2_X1 g_g5564 (I10018, I10019, g5564);
NAND2_X1 g_g5565 (g2044, g4933, g5565);
NAND2_X1 g_g5567 (g1879, g4883, g5567);
NAND3_X1 g_g5568 (g2044, g4902, g4320, g5568);
NAND2_X1 g_I10038 (g4893, g2202, I10038);
NAND2_X1 g_I10039 (g4893, I10038, I10039);
NAND2_X1 g_I10040 (g2202, I10038, I10040);
NAND2_X1 g_g5575 (I10039, I10040, g5575);
NAND3_X1 g_g5576 (g4894, g4888, g4884, g5576);
NAND2_X1 g_I10060 (g4910, g2226, I10060);
NAND2_X1 g_I10061 (g4910, I10060, I10061);
NAND2_X1 g_I10062 (g2226, I10060, I10062);
NAND2_X1 g_g5589 (I10061, I10062, g5589);
NAND2_X1 g_g5590 (g2044, g4906, g5590);
NAND2_X1 g_I10071 (g4954, g2253, I10071);
NAND2_X1 g_I10072 (g4954, I10071, I10072);
NAND2_X1 g_I10073 (g2253, I10071, I10073);
NAND2_X1 g_g5594 (I10072, I10073, g5594);
NAND2_X1 g_I10078 (g4911, g2256, I10078);
NAND2_X1 g_I10079 (g4911, I10078, I10079);
NAND2_X1 g_I10080 (g2256, I10078, I10080);
NAND2_X1 g_g5595 (I10079, I10080, g5595);
NAND2_X1 g_I10092 (g4881, g2177, I10092);
NAND2_X1 g_I10093 (g4881, I10092, I10093);
NAND2_X1 g_I10094 (g2177, I10092, I10094);
NAND2_X1 g_g5605 (I10093, I10094, g5605);
NAND2_X1 g_g5625 (g2044, g4957, g5625);
NAND2_X1 g_g5632 (g2276, g4901, g5632);
NAND2_X1 g_g5657 (g5021, g4381, g5657);
NAND2_X1 g_I10142 (g4707, g1916, I10142);
NAND2_X1 g_I10143 (g4707, I10142, I10143);
NAND2_X1 g_I10144 (g1916, I10142, I10144);
NAND2_X1 g_g5661 (I10143, I10144, g5661);
NAND3_X1 g_g5672 (g5056, g5039, g5023, g5672);
NAND2_X1 g_g5681 (g5132, g2043, g5681);
NAND2_X1 g_g5686 (g5132, g1263, g5686);
NAND2_X1 g_I10196 (g4724, g1958, I10196);
NAND2_X1 g_I10197 (g4724, I10196, I10197);
NAND2_X1 g_I10198 (g1958, I10196, I10198);
NAND2_X1 g_g5689 (I10197, I10198, g5689);
NAND2_X1 g_g5697 (g2044, g5005, g5697);
NAND2_X1 g_I10223 (g2522, g4895, I10223);
NAND2_X1 g_I10224 (g2522, I10223, I10224);
NAND2_X1 g_I10225 (g4895, I10223, I10225);
NAND2_X1 g_g5712 (I10224, I10225, g5712);
NAND2_X1 g_I10298 (g5461, g2562, I10298);
NAND2_X1 g_I10299 (g5461, I10298, I10299);
NAND2_X1 g_I10300 (g2562, I10298, I10300);
NAND2_X1 g_g5747 (I10299, I10300, g5747);
NAND2_X1 g_I10305 (g5470, g3019, I10305);
NAND2_X1 g_I10306 (g5470, I10305, I10306);
NAND2_X1 g_I10307 (g3019, I10305, I10307);
NAND2_X1 g_g5748 (I10306, I10307, g5748);
NAND2_X1 g_I10313 (g5484, g1041, I10313);
NAND2_X1 g_I10314 (g5484, I10313, I10314);
NAND2_X1 g_I10315 (g1041, I10313, I10315);
NAND2_X1 g_g5750 (I10314, I10315, g5750);
NAND2_X1 g_I10320 (g5459, g2573, I10320);
NAND2_X1 g_I10321 (g5459, I10320, I10321);
NAND2_X1 g_I10322 (g2573, I10320, I10322);
NAND2_X1 g_g5751 (I10321, I10322, g5751);
NAND2_X1 g_I10327 (g5467, g2562, I10327);
NAND2_X1 g_I10328 (g5467, I10327, I10328);
NAND2_X1 g_I10329 (g2562, I10327, I10329);
NAND2_X1 g_g5752 (I10328, I10329, g5752);
NAND2_X1 g_I10334 (g5462, g2573, I10334);
NAND2_X1 g_I10335 (g5462, I10334, I10335);
NAND2_X1 g_I10336 (g2573, I10334, I10336);
NAND2_X1 g_g5753 (I10335, I10336, g5753);
NAND2_X1 g_I10359 (g5552, g1118, I10359);
NAND2_X1 g_I10360 (g5552, I10359, I10360);
NAND2_X1 g_I10361 (g1118, I10359, I10361);
NAND2_X1 g_g5762 (I10360, I10361, g5762);
NAND2_X1 g_I10625 (g5314, g1514, I10625);
NAND2_X1 g_I10626 (g5314, I10625, I10626);
NAND2_X1 g_I10627 (g1514, I10625, I10627);
NAND2_X1 g_g6023 (I10626, I10627, g6023);
NAND2_X1 g_I10743 (g5550, g2100, I10743);
NAND2_X1 g_I10744 (g5550, I10743, I10744);
NAND2_X1 g_I10745 (g2100, I10743, I10745);
NAND2_X1 g_g6119 (I10744, I10745, g6119);
NAND2_X1 g_I10789 (g5512, g2170, I10789);
NAND2_X1 g_I10790 (g5512, I10789, I10790);
NAND2_X1 g_I10791 (g2170, I10789, I10791);
NAND2_X1 g_g6142 (I10790, I10791, g6142);
NAND2_X1 g_I10818 (g5567, g2039, I10818);
NAND2_X1 g_I10819 (g5567, I10818, I10819);
NAND2_X1 g_I10820 (g2039, I10818, I10820);
NAND2_X1 g_g6153 (I10819, I10820, g6153);
NAND4_X1 g_g6158 (g3735, g3716, g5633, g3754, g6158);
NAND2_X1 g_I10834 (g5514, g2584, I10834);
NAND2_X1 g_I10835 (g5514, I10834, I10835);
NAND2_X1 g_I10836 (g2584, I10834, I10836);
NAND2_X1 g_g6159 (I10835, I10836, g6159);
NAND2_X1 g_g6163 (g5633, g3716, g6163);
NAND2_X1 g_I10847 (g5490, g2595, I10847);
NAND2_X1 g_I10848 (g5490, I10847, I10848);
NAND2_X1 g_I10849 (g2595, I10847, I10849);
NAND2_X1 g_g6164 (I10848, I10849, g6164);
NAND2_X1 g_I10854 (g5521, g2584, I10854);
NAND2_X1 g_I10855 (g5521, I10854, I10855);
NAND2_X1 g_I10856 (g2584, I10854, I10856);
NAND2_X1 g_g6165 (I10855, I10856, g6165);
NAND2_X1 g_I10866 (g5480, g2605, I10866);
NAND2_X1 g_I10867 (g5480, I10866, I10867);
NAND2_X1 g_I10868 (g2605, I10866, I10868);
NAND2_X1 g_g6169 (I10867, I10868, g6169);
NAND2_X1 g_I10873 (g5516, g2595, I10873);
NAND2_X1 g_I10874 (g5516, I10873, I10874);
NAND2_X1 g_I10875 (g2595, I10873, I10875);
NAND2_X1 g_g6170 (I10874, I10875, g6170);
NAND2_X1 g_I10888 (g5590, g2259, I10888);
NAND2_X1 g_I10889 (g5590, I10888, I10889);
NAND2_X1 g_I10890 (g2259, I10888, I10890);
NAND2_X1 g_g6177 (I10889, I10890, g6177);
NAND2_X1 g_g6178 (g2205, g5568, g6178);
NAND2_X1 g_I10899 (g5520, g2752, I10899);
NAND2_X1 g_I10900 (g5520, I10899, I10900);
NAND2_X1 g_I10901 (g2752, I10899, I10901);
NAND2_X1 g_g6180 (I10900, I10901, g6180);
NAND2_X1 g_I10906 (g5492, g2605, I10906);
NAND2_X1 g_I10907 (g5492, I10906, I10907);
NAND2_X1 g_I10908 (g2605, I10906, I10908);
NAND2_X1 g_g6181 (I10907, I10908, g6181);
NAND3_X1 g_g6187 (g5633, g3735, g3716, g6187);
NAND2_X1 g_I10923 (g5525, g2752, I10923);
NAND2_X1 g_I10924 (g5525, I10923, I10924);
NAND2_X1 g_I10925 (g2752, I10923, I10925);
NAND2_X1 g_g6188 (I10924, I10925, g6188);
NAND2_X1 g_I10952 (g5565, g2340, I10952);
NAND2_X1 g_I10953 (g5565, I10952, I10953);
NAND2_X1 g_I10954 (g2340, I10952, I10954);
NAND2_X1 g_g6203 (I10953, I10954, g6203);
NAND2_X1 g_I10980 (g5625, g2210, I10980);
NAND2_X1 g_I10981 (g5625, I10980, I10981);
NAND2_X1 g_I10982 (g2210, I10980, I10982);
NAND2_X1 g_g6215 (I10981, I10982, g6215);
NAND2_X1 g_I10991 (g5632, g2389, I10991);
NAND2_X1 g_I10992 (g5632, I10991, I10992);
NAND2_X1 g_I10993 (g2389, I10991, I10993);
NAND2_X1 g_g6218 (I10992, I10993, g6218);
NAND2_X1 g_I11078 (g5697, g2511, I11078);
NAND2_X1 g_I11079 (g5697, I11078, I11079);
NAND2_X1 g_I11080 (g2511, I11078, I11080);
NAND2_X1 g_g6265 (I11079, I11080, g6265);
NAND2_X1 g_I11094 (g5515, g2734, I11094);
NAND2_X1 g_I11095 (g5515, I11094, I11095);
NAND2_X1 g_I11096 (g2734, I11094, I11096);
NAND2_X1 g_g6273 (I11095, I11096, g6273);
NAND2_X1 g_I11101 (g5491, g2712, I11101);
NAND2_X1 g_I11102 (g5491, I11101, I11102);
NAND2_X1 g_I11103 (g2712, I11101, I11103);
NAND2_X1 g_g6274 (I11102, I11103, g6274);
NAND2_X1 g_I11108 (g5522, g2734, I11108);
NAND2_X1 g_I11109 (g5522, I11108, I11109);
NAND2_X1 g_I11110 (g2734, I11108, I11110);
NAND2_X1 g_g6275 (I11109, I11110, g6275);
NAND2_X1 g_I11115 (g5481, g3062, I11115);
NAND2_X1 g_I11116 (g5481, I11115, I11116);
NAND2_X1 g_I11117 (g3062, I11115, I11117);
NAND2_X1 g_g6276 (I11116, I11117, g6276);
NAND2_X1 g_I11122 (g5517, g2712, I11122);
NAND2_X1 g_I11123 (g5517, I11122, I11123);
NAND2_X1 g_I11124 (g2712, I11122, I11124);
NAND2_X1 g_g6277 (I11123, I11124, g6277);
NAND2_X1 g_I11135 (g5476, g3052, I11135);
NAND2_X1 g_I11136 (g5476, I11135, I11136);
NAND2_X1 g_I11137 (g3052, I11135, I11137);
NAND2_X1 g_g6280 (I11136, I11137, g6280);
NAND2_X1 g_I11142 (g5493, g3062, I11142);
NAND2_X1 g_I11143 (g5493, I11142, I11143);
NAND2_X1 g_I11144 (g3062, I11142, I11144);
NAND2_X1 g_g6281 (I11143, I11144, g6281);
NAND2_X1 g_I11149 (g5473, g3038, I11149);
NAND2_X1 g_I11150 (g5473, I11149, I11150);
NAND2_X1 g_I11151 (g3038, I11149, I11151);
NAND2_X1 g_g6282 (I11150, I11151, g6282);
NAND2_X1 g_I11156 (g5482, g3052, I11156);
NAND2_X1 g_I11157 (g5482, I11156, I11157);
NAND2_X1 g_I11158 (g3052, I11156, I11158);
NAND2_X1 g_g6283 (I11157, I11158, g6283);
NAND2_X1 g_I11163 (g5469, g3029, I11163);
NAND2_X1 g_I11164 (g5469, I11163, I11164);
NAND2_X1 g_I11165 (g3029, I11163, I11165);
NAND2_X1 g_g6284 (I11164, I11165, g6284);
NAND2_X1 g_I11170 (g5477, g3038, I11170);
NAND2_X1 g_I11171 (g5477, I11170, I11171);
NAND2_X1 g_I11172 (g3038, I11170, I11172);
NAND2_X1 g_g6285 (I11171, I11172, g6285);
NAND2_X1 g_I11177 (g5466, g3019, I11177);
NAND2_X1 g_I11178 (g5466, I11177, I11178);
NAND2_X1 g_I11179 (g3019, I11177, I11179);
NAND2_X1 g_g6286 (I11178, I11179, g6286);
NAND2_X1 g_I11184 (g5474, g3029, I11184);
NAND2_X1 g_I11185 (g5474, I11184, I11185);
NAND2_X1 g_I11186 (g3029, I11184, I11186);
NAND2_X1 g_g6287 (I11185, I11186, g6287);
NAND2_X1 g_I11549 (g5984, g1045, I11549);
NAND2_X1 g_I11550 (g5984, I11549, I11550);
NAND2_X1 g_I11551 (g1045, I11549, I11551);
NAND2_X1 g_g6424 (I11550, I11551, g6424);
NAND2_X1 g_I11574 (g5894, g1122, I11574);
NAND2_X1 g_I11575 (g5894, I11574, I11575);
NAND2_X1 g_I11576 (g1122, I11574, I11576);
NAND2_X1 g_g6435 (I11575, I11576, g6435);
NAND2_X1 g_g6463 (g5918, g5278, g6463);
NAND2_X1 g_I11614 (g6239, g1519, I11614);
NAND2_X1 g_I11615 (g6239, I11614, I11615);
NAND2_X1 g_I11616 (g1519, I11614, I11616);
NAND2_X1 g_g6466 (I11615, I11616, g6466);
NAND2_X1 g_g6467 (g5956, g5269, g6467);
NAND2_X1 g_g6469 (g5918, g5278, g6469);
NAND2_X1 g_g6472 (g5971, g5269, g6472);
NAND2_X1 g_g6473 (g5269, g5988, g6473);
NAND2_X1 g_g6476 (g5939, g5269, g6476);
NAND2_X1 g_g6477 (g5269, g5918, g6477);
NAND2_X1 g_g6482 (g5269, g5847, g6482);
NAND2_X1 g_g6497 (g5278, g5847, g6497);
NAND2_X1 g_g6503 (g5269, g5897, g6503);
NAND2_X1 g_g6504 (g5269, g5874, g6504);
NAND2_X1 g_g6510 (g5278, g5874, g6510);
NAND2_X1 g_g6516 (g5897, g5278, g6516);
NAND2_X1 g_g6559 (g5814, g6109, g6559);
NAND2_X1 g_I11750 (g6112, g1486, I11750);
NAND2_X1 g_I11751 (g6112, I11750, I11751);
NAND2_X1 g_I11752 (g1486, I11750, I11752);
NAND2_X1 g_g6570 (I11751, I11752, g6570);
NAND2_X1 g_I11757 (g1758, g6118, I11757);
NAND2_X1 g_I11758 (g1758, I11757, I11758);
NAND2_X1 g_I11759 (g6118, I11757, I11759);
NAND2_X1 g_g6571 (I11758, I11759, g6571);
NAND2_X1 g_I11841 (g2548, g6158, I11841);
NAND2_X1 g_I11842 (g2548, I11841, I11842);
NAND2_X1 g_I11843 (g6158, I11841, I11843);
NAND2_X1 g_g6615 (I11842, I11843, g6615);
NAND2_X1 g_I11873 (g2543, g6187, I11873);
NAND2_X1 g_I11874 (g2543, I11873, I11874);
NAND2_X1 g_I11875 (g6187, I11873, I11875);
NAND2_X1 g_g6627 (I11874, I11875, g6627);
NAND2_X1 g_g6680 (g5403, g6252, g6680);
NAND2_X1 g_I12015 (g5874, g5847, I12015);
NAND2_X1 g_I12016 (g5874, I12015, I12016);
NAND2_X1 g_I12017 (g5847, I12015, I12017);
NAND2_X1 g_g6695 (I12016, I12017, g6695);
NAND2_X1 g_I12031 (g5918, g5897, I12031);
NAND2_X1 g_I12032 (g5918, I12031, I12032);
NAND2_X1 g_I12033 (g5897, I12031, I12033);
NAND2_X1 g_g6701 (I12032, I12033, g6701);
NAND2_X1 g_I12051 (g5956, g5939, I12051);
NAND2_X1 g_I12052 (g5956, I12051, I12052);
NAND2_X1 g_I12053 (g5939, I12051, I12053);
NAND2_X1 g_g6709 (I12052, I12053, g6709);
NAND2_X1 g_I12078 (g5988, g5971, I12078);
NAND2_X1 g_I12079 (g5988, I12078, I12079);
NAND2_X1 g_I12080 (g5971, I12078, I12080);
NAND2_X1 g_g6722 (I12079, I12080, g6722);
NAND2_X1 g_I12179 (g1961, g6163, I12179);
NAND2_X1 g_I12180 (g1961, I12179, I12180);
NAND2_X1 g_I12181 (g6163, I12179, I12181);
NAND2_X1 g_g6770 (I12180, I12181, g6770);
NAND2_X1 g_I12550 (g6689, g1462, I12550);
NAND2_X1 g_I12551 (g6689, I12550, I12551);
NAND2_X1 g_I12552 (g1462, I12550, I12552);
NAND2_X1 g_g6893 (I12551, I12552, g6893);
NAND2_X1 g_I12575 (g6574, g1049, I12575);
NAND2_X1 g_I12576 (g6574, I12575, I12576);
NAND2_X1 g_I12577 (g1049, I12575, I12577);
NAND2_X1 g_g6902 (I12576, I12577, g6902);
NAND2_X1 g_I12596 (g6582, g1126, I12596);
NAND2_X1 g_I12597 (g6582, I12596, I12597);
NAND2_X1 g_I12598 (g1126, I12596, I12598);
NAND2_X1 g_g6911 (I12597, I12598, g6911);
NAND2_X1 g_I12832 (g6722, g6709, I12832);
NAND2_X1 g_I12833 (g6722, I12832, I12833);
NAND2_X1 g_I12834 (g6709, I12832, I12834);
NAND2_X1 g_g7065 (I12833, I12834, g7065);
NAND2_X1 g_g7069 (g5435, g6680, g7069);
NAND2_X1 g_I12852 (g6701, g6695, I12852);
NAND2_X1 g_I12853 (g6701, I12852, I12853);
NAND2_X1 g_I12854 (g6695, I12852, I12854);
NAND2_X1 g_g7082 (I12853, I12854, g7082);
NAND2_X1 g_I12869 (g2536, g6618, I12869);
NAND2_X1 g_I12870 (g2536, I12869, I12870);
NAND2_X1 g_I12871 (g6618, I12869, I12871);
NAND2_X1 g_g7093 (I12870, I12871, g7093);
NAND2_X1 g_I12951 (g7003, g1467, I12951);
NAND2_X1 g_I12952 (g7003, I12951, I12952);
NAND2_X1 g_I12953 (g1467, I12951, I12953);
NAND2_X1 g_g7121 (I12952, I12953, g7121);
NAND2_X1 g_I13002 (g7010, g1053, I13002);
NAND2_X1 g_I13003 (g7010, I13002, I13003);
NAND2_X1 g_I13004 (g1053, I13002, I13004);
NAND2_X1 g_g7140 (I13003, I13004, g7140);
NAND2_X1 g_I13016 (g6941, g1142, I13016);
NAND2_X1 g_I13017 (g6941, I13016, I13017);
NAND2_X1 g_I13018 (g1142, I13016, I13018);
NAND2_X1 g_g7144 (I13017, I13018, g7144);
NAND4_X1 g_g7234 (g3757, g3739, g7050, g3770, g7234);
NAND2_X1 g_g7237 (g7050, g3739, g7237);
NAND3_X1 g_g7244 (g7050, g3757, g3739, g7244);
NAND2_X1 g_I13213 (g7065, g7082, I13213);
NAND2_X1 g_I13214 (g7065, I13213, I13214);
NAND2_X1 g_I13215 (g7082, I13213, I13215);
NAND2_X1 g_g7257 (I13214, I13215, g7257);
NAND2_X1 g_I13376 (g7199, g1472, I13376);
NAND2_X1 g_I13377 (g7199, I13376, I13377);
NAND2_X1 g_I13378 (g1472, I13376, I13378);
NAND2_X1 g_g7316 (I13377, I13378, g7316);
NAND2_X1 g_I13395 (g7212, g1057, I13395);
NAND2_X1 g_I13396 (g7212, I13395, I13396);
NAND2_X1 g_I13397 (g1057, I13395, I13397);
NAND2_X1 g_g7325 (I13396, I13397, g7325);
NAND2_X1 g_I13587 (g2556, g7234, I13587);
NAND2_X1 g_I13588 (g2556, I13587, I13588);
NAND2_X1 g_I13589 (g7234, I13587, I13589);
NAND2_X1 g_g7444 (I13588, I13589, g7444);
NAND2_X1 g_I13598 (g2551, g7244, I13598);
NAND2_X1 g_I13599 (g2551, I13598, I13599);
NAND2_X1 g_I13600 (g7244, I13598, I13600);
NAND2_X1 g_g7447 (I13599, I13600, g7447);
NAND2_X1 g_I13638 (g7257, g7069, I13638);
NAND2_X1 g_I13639 (g7257, I13638, I13639);
NAND2_X1 g_I13640 (g7069, I13638, I13640);
NAND2_X1 g_g7480 (I13639, I13640, g7480);
NAND2_X1 g_I13685 (g1977, g7237, I13685);
NAND2_X1 g_I13686 (g1977, I13685, I13686);
NAND2_X1 g_I13687 (g7237, I13685, I13687);
NAND2_X1 g_g7503 (I13686, I13687, g7503);
NAND2_X1 g_I13785 (g7427, g1477, I13785);
NAND2_X1 g_I13786 (g7427, I13785, I13786);
NAND2_X1 g_I13787 (g1477, I13785, I13787);
NAND2_X1 g_g7535 (I13786, I13787, g7535);
NAND2_X1 g_I13800 (g7429, g1061, I13800);
NAND2_X1 g_I13801 (g7429, I13800, I13801);
NAND2_X1 g_I13802 (g1061, I13800, I13802);
NAND2_X1 g_g7540 (I13801, I13802, g7540);
NAND2_X1 g_I14244 (g7683, g1065, I14244);
NAND2_X1 g_I14245 (g7683, I14244, I14245);
NAND2_X1 g_I14246 (g1065, I14244, I14246);
NAND2_X1 g_g7828 (I14245, I14246, g7828);
NAND2_X1 g_I14472 (g8147, g1069, I14472);
NAND2_X1 g_I14473 (g8147, I14472, I14473);
NAND2_X1 g_I14474 (g1069, I14472, I14474);
NAND2_X1 g_g8231 (I14473, I14474, g8231);
NAND2_X1 g_g8239 (g8073, g8092, g8239);
NAND2_X1 g_g8627 (g6232, g8091, g8627);
NAND2_X1 g_g8633 (g8176, g6232, g8633);
NAND2_X1 g_I14837 (g8660, g1073, I14837);
NAND2_X1 g_I14838 (g8660, I14837, I14838);
NAND2_X1 g_I14839 (g1073, I14837, I14839);
NAND2_X1 g_g8681 (I14838, I14839, g8681);
NAND2_X1 g_g8798 (g6984, g8644, g8798);
NAND2_X1 g_I15817 (g9151, g9148, I15817);
NAND2_X1 g_I15818 (g9151, I15817, I15818);
NAND2_X1 g_I15819 (g9148, I15817, I15819);
NAND2_X1 g_g9179 (I15818, I15819, g9179);
NAND2_X1 g_I15848 (g9162, g9154, I15848);
NAND2_X1 g_I15849 (g9162, I15848, I15849);
NAND2_X1 g_I15850 (g9154, I15848, I15850);
NAND2_X1 g_g9190 (I15849, I15850, g9190);
NAND2_X1 g_I15855 (g9168, g9165, I15855);
NAND2_X1 g_I15856 (g9168, I15855, I15856);
NAND2_X1 g_I15857 (g9165, I15855, I15857);
NAND2_X1 g_g9191 (I15856, I15857, g9191);
NAND2_X1 g_I15862 (g9174, g9171, I15862);
NAND2_X1 g_I15863 (g9174, I15862, I15863);
NAND2_X1 g_I15864 (g9171, I15862, I15864);
NAND2_X1 g_g9192 (I15863, I15864, g9192);
NAND2_X1 g_I15880 (g9190, g9179, I15880);
NAND2_X1 g_I15881 (g9190, I15880, I15881);
NAND2_X1 g_I15882 (g9179, I15880, I15882);
NAND2_X1 g_g9202 (I15881, I15882, g9202);
NAND2_X1 g_I15887 (g9192, g9191, I15887);
NAND2_X1 g_I15888 (g9192, I15887, I15888);
NAND2_X1 g_I15889 (g9191, I15887, I15889);
NAND2_X1 g_g9203 (I15888, I15889, g9203);
NAND2_X1 g_I15897 (g9202, g9203, I15897);
NAND2_X1 g_I15898 (g9202, I15897, I15898);
NAND2_X1 g_I15899 (g9203, I15897, I15899);
NAND2_X1 g_g9205 (I15898, I15899, g9205);
NOR2_X1 g_g1964 (g1428, g1429, g1964);
NOR2_X1 g_g1980 (g1430, g1431, g1980);
NOR2_X1 g_g2014 (g1421, g1416, g2014);
NOR2_X1 g_g2521 (g65, g62, g2521);
NOR3_X1 g_g3225 (g1021, g1025, g1889, g3225);
NOR2_X1 g_g3233 (g1714, g1459, g3233);
NOR3_X1 g_g3237 (g1444, g1838, g1454, g3237);
NOR2_X1 g_g3260 (g1728, g2490, g3260);
NOR2_X1 g_g3310 (g936, g2557, g3310);
NOR4_X1 g_g3504 (g1375, g2229, g2213, g2206, g3504);
NOR2_X1 g_g3505 (g2263, g1395, g3505);
NOR4_X1 g_g3515 (g1388, g2262, g2230, g2214, g3515);
NOR2_X1 g_g3516 (g2282, g1401, g3516);
NOR2_X1 g_g3528 (g2343, g1391, g3528);
NOR2_X1 g_g3555 (g2359, g1398, g3555);
NOR3_X1 g_g3790 (g985, g990, g2295, g3790);
NOR2_X1 g_g3885 (g3310, g3466, g3885);
NOR2_X1 g_g4160 (g1231, g2834, g4160);
NOR2_X1 g_g4232 (g1934, g3591, g4232);
NOR2_X1 g_g4318 (g3681, g1590, g4318);
NOR2_X1 g_g4349 (g2496, g3310, g4349);
NOR2_X1 g_g4354 (g1424, g3541, g4354);
NOR2_X1 g_g4676 (g3885, g3094, g4676);
NOR4_X1 g_g4884 (g4492, g4476, g4456, g4294, g4884);
NOR4_X1 g_g4888 (g4548, g4528, g4513, g4502, g4888);
NOR3_X1 g_g4894 (g4298, g4575, g4563, g4894);
NOR4_X1 g_g5023 (g3894, g3889, g3886, g4359, g5023);
NOR4_X1 g_g5039 (g3924, g3914, g3906, g3899, g5039);
NOR3_X1 g_g5056 (g3556, g2872, g3938, g5056);
NOR3_X1 g_g5614 (g3002, g1590, g4714, g5614);
NOR2_X1 g_g5615 (g4714, g3002, g5615);
NOR2_X1 g_g5772 (g5428, g1888, g5772);
NOR2_X1 g_g6174 (g1855, g5305, g6174);
NOR2_X1 g_g6184 (g875, g5291, g6184);
NOR2_X1 g_g6185 (g5305, g1590, g6185);
NOR2_X1 g_g6193 (g1926, g5310, g6193);
NOR4_X1 g_g6197 (g875, g866, g1590, g5291, g6197);
NOR2_X1 g_g6209 (g2332, g5305, g6209);
NOR2_X1 g_g6214 (g878, g5284, g6214);
NOR2_X1 g_g6259 (g3002, g5312, g6259);
NOR2_X1 g_g6452 (g6270, g2245, g6452);
NOR4_X1 g_g6465 (g5403, g5802, g5769, g5790, g6465);
NOR3_X1 g_g6489 (g5802, g5769, g5790, g6489);
NOR3_X1 g_g6664 (g5836, g1901, g1788, g6664);
NOR4_X1 g_g6910 (g1011, g1837, g6559, g1008, g6910);
NOR3_X1 g_g7152 (g6253, g7083, g5418, g7152);
NOR3_X1 g_g7209 (g1789, g146, g6984, g7209);
NOR2_X1 g_g7312 (g7178, g6970, g7312);
NOR2_X1 g_g7314 (g7180, g6972, g7314);
NOR2_X1 g_g7318 (g7185, g6979, g7318);
NOR2_X1 g_g7321 (g7187, g6990, g7321);
NOR2_X1 g_g7322 (g7188, g6991, g7322);
NOR2_X1 g_g7324 (g7189, g6994, g7324);
NOR2_X1 g_g7326 (g7194, g6999, g7326);
NOR2_X1 g_g7328 (g7196, g7001, g7328);
NOR2_X1 g_g7406 (g7191, g1600, g7406);
NOR2_X1 g_g7566 (g7421, g1597, g7566);
NOR2_X1 g_g8073 (g7658, g7654, g8073);
NOR4_X1 g_g8092 (g7634, g7628, g7616, g7611, g8092);
NOR3_X1 g_g8230 (g8199, I14467, I14468, g8230);
NOR3_X1 g_g8232 (g8199, I14479, I14480, g8232);
NOR3_X1 g_g8233 (g8199, I14484, I14485, g8233);
NOR3_X1 g_g8236 (g8199, I14495, I14496, g8236);
NOR4_X1 g_g8279 (g7658, g7616, g8082, g7634, g8279);
NOR4_X1 g_g8360 (g7658, g7616, g8082, g7634, g8360);
NOR4_X1 g_g8523 (g7658, g7616, g8082, g7634, g8523);
NOR4_X1 g_g8625 (g1000, g6573, g1860, g8009, g8625);
NOR2_X1 g_g8629 (g6270, g8009, g8629);
NOR4_X1 g_g8630 (g6110, g7784, g3591, g1864, g8630);
NOR2_X1 g_g8635 (g1034, g8128, g8635);
NOR4_X1 g_g8641 (g6559, g162, g7784, g3591, g8641);
NOR2_X1 g_g8644 (g4146, g8128, g8644);
NOR3_X1 g_g8655 (g8199, I14753, I14754, g8655);
NOR3_X1 g_g8656 (g8199, I14758, I14759, g8656);
NOR3_X1 g_g8658 (g8199, I14766, I14767, g8658);
NOR3_X1 g_g8659 (g8199, I14771, I14772, g8659);
NOR3_X1 g_g8679 (g8493, g8239, I14831, g8679);
NOR3_X1 g_g8680 (g8493, g8239, I14834, g8680);
NOR3_X1 g_g8694 (g7658, g8613, g7634, g8694);
NOR3_X1 g_g8699 (g7658, g8613, g7634, g8699);
NOR3_X1 g_g8706 (g7658, g8613, g7634, g8706);
NOR3_X1 g_g8707 (g7658, g8613, g7634, g8707);
NOR2_X1 g_g8801 (g8635, g3790, g8801);
NOR3_X1 g_g8803 (g8443, g8421, I15021, g8803);
NOR3_X1 g_g8805 (g8443, g8421, I15033, g8805);
NOR3_X1 g_g8806 (g8443, g8421, I15044, g8806);
NOR3_X1 g_g8807 (g8443, g8421, I15055, g8807);
NOR3_X1 g_g8811 (g8443, g8421, I15075, g8811);
NOR3_X1 g_g8812 (g8443, g8421, I15086, g8812);
NOR3_X1 g_g8818 (g8443, g8421, I15102, g8818);
NOR3_X1 g_g8819 (g8443, g8421, I15113, g8819);
NOR3_X1 g_g8847 (g8493, g8239, I15147, g8847);
NOR3_X1 g_g8850 (g8493, g8239, I15152, g8850);
NOR3_X1 g_g8855 (g7658, g8613, g7634, g8855);
NOR3_X1 g_g8859 (g8493, g8239, I15165, g8859);
NOR3_X1 g_g8861 (g8493, g8239, I15169, g8861);
NOR3_X1 g_g8862 (g8493, g8239, I15172, g8862);
NOR3_X1 g_g8863 (g8493, g8239, I15175, g8863);
endmodule
